
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_MUX21_GENERIC_N16_1 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_MUX21_GENERIC_N16_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_47 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_47;

architecture SYN_behavioral of NAND2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_46 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_46;

architecture SYN_behavioral of NAND2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_45 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_45;

architecture SYN_behavioral of NAND2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_44 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_44;

architecture SYN_behavioral of NAND2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_43 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_43;

architecture SYN_behavioral of NAND2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_42 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_42;

architecture SYN_behavioral of NAND2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_41 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_41;

architecture SYN_behavioral of NAND2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_40 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_40;

architecture SYN_behavioral of NAND2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_39 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_39;

architecture SYN_behavioral of NAND2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_38 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_38;

architecture SYN_behavioral of NAND2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_37 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_37;

architecture SYN_behavioral of NAND2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_36 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_36;

architecture SYN_behavioral of NAND2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_35 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_35;

architecture SYN_behavioral of NAND2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_34 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_34;

architecture SYN_behavioral of NAND2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_33 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_33;

architecture SYN_behavioral of NAND2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_32 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_32;

architecture SYN_behavioral of NAND2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_31 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_31;

architecture SYN_behavioral of NAND2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_30 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_30;

architecture SYN_behavioral of NAND2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_29 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_29;

architecture SYN_behavioral of NAND2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_28 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_28;

architecture SYN_behavioral of NAND2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_27 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_27;

architecture SYN_behavioral of NAND2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_26 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_26;

architecture SYN_behavioral of NAND2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_25 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_25;

architecture SYN_behavioral of NAND2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_24 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_24;

architecture SYN_behavioral of NAND2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_23 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_23;

architecture SYN_behavioral of NAND2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_22 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_22;

architecture SYN_behavioral of NAND2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_21 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_21;

architecture SYN_behavioral of NAND2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_20 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_20;

architecture SYN_behavioral of NAND2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_19 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_19;

architecture SYN_behavioral of NAND2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_18 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_18;

architecture SYN_behavioral of NAND2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_17 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_17;

architecture SYN_behavioral of NAND2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_16 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_16;

architecture SYN_behavioral of NAND2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_15 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_15;

architecture SYN_behavioral of NAND2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_14 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_14;

architecture SYN_behavioral of NAND2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_13 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_13;

architecture SYN_behavioral of NAND2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_12 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_12;

architecture SYN_behavioral of NAND2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_11 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_11;

architecture SYN_behavioral of NAND2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_10 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_10;

architecture SYN_behavioral of NAND2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_9 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_9;

architecture SYN_behavioral of NAND2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_8 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_8;

architecture SYN_behavioral of NAND2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_7 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_7;

architecture SYN_behavioral of NAND2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_6 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_6;

architecture SYN_behavioral of NAND2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_5 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_5;

architecture SYN_behavioral of NAND2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_4 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_4;

architecture SYN_behavioral of NAND2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_3 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_3;

architecture SYN_behavioral of NAND2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_2 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_2;

architecture SYN_behavioral of NAND2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_1 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_1;

architecture SYN_behavioral of NAND2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity NAND2_0 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_0;

architecture SYN_behavioral of NAND2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity INV is

   port( a : in std_logic;  f : out std_logic);

end INV;

architecture SYN_behavioral of INV is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X1 port map( A => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_MUX21_GENERIC_N16_1.all;

entity MUX21_GENERIC_N16_1 is

   port( A, B : in std_logic_vector (15 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (15 downto 0));

end MUX21_GENERIC_N16_1;

architecture SYN_structural of MUX21_GENERIC_N16_1 is

   component NAND2_1
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_2
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_3
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_4
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_5
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_6
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_7
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_8
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_9
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_10
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_11
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_12
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_13
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_14
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_15
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_16
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_17
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_18
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_19
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_20
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_21
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_22
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_23
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_24
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_25
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_26
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_27
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_28
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_29
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_30
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_31
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_32
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_33
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_34
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_35
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_36
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_37
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_38
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_39
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_40
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_41
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_42
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_43
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_44
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_45
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_46
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_47
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_0
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component INV
      port( a : in std_logic;  f : out std_logic);
   end component;
   
   signal sel_not, s1_15_port, s1_14_port, s1_13_port, s1_12_port, s1_11_port, 
      s1_10_port, s1_9_port, s1_8_port, s1_7_port, s1_6_port, s1_5_port, 
      s1_4_port, s1_3_port, s1_2_port, s1_1_port, s1_0_port, s2_15_port, 
      s2_14_port, s2_13_port, s2_12_port, s2_11_port, s2_10_port, s2_9_port, 
      s2_8_port, s2_7_port, s2_6_port, s2_5_port, s2_4_port, s2_3_port, 
      s2_2_port, s2_1_port, s2_0_port : std_logic;

begin
   
   inv_sel : INV port map( a => SEL, f => sel_not);
   s1_i_0 : NAND2_0 port map( a => A(0), b => sel_not, f => s1_0_port);
   s2_i_0 : NAND2_47 port map( a => B(0), b => SEL, f => s2_0_port);
   y_i_0 : NAND2_46 port map( a => s1_0_port, b => s2_0_port, f => Y(0));
   s1_i_1 : NAND2_45 port map( a => A(1), b => sel_not, f => s1_1_port);
   s2_i_1 : NAND2_44 port map( a => B(1), b => SEL, f => s2_1_port);
   y_i_1 : NAND2_43 port map( a => s1_1_port, b => s2_1_port, f => Y(1));
   s1_i_2 : NAND2_42 port map( a => A(2), b => sel_not, f => s1_2_port);
   s2_i_2 : NAND2_41 port map( a => B(2), b => SEL, f => s2_2_port);
   y_i_2 : NAND2_40 port map( a => s1_2_port, b => s2_2_port, f => Y(2));
   s1_i_3 : NAND2_39 port map( a => A(3), b => sel_not, f => s1_3_port);
   s2_i_3 : NAND2_38 port map( a => B(3), b => SEL, f => s2_3_port);
   y_i_3 : NAND2_37 port map( a => s1_3_port, b => s2_3_port, f => Y(3));
   s1_i_4 : NAND2_36 port map( a => A(4), b => sel_not, f => s1_4_port);
   s2_i_4 : NAND2_35 port map( a => B(4), b => SEL, f => s2_4_port);
   y_i_4 : NAND2_34 port map( a => s1_4_port, b => s2_4_port, f => Y(4));
   s1_i_5 : NAND2_33 port map( a => A(5), b => sel_not, f => s1_5_port);
   s2_i_5 : NAND2_32 port map( a => B(5), b => SEL, f => s2_5_port);
   y_i_5 : NAND2_31 port map( a => s1_5_port, b => s2_5_port, f => Y(5));
   s1_i_6 : NAND2_30 port map( a => A(6), b => sel_not, f => s1_6_port);
   s2_i_6 : NAND2_29 port map( a => B(6), b => SEL, f => s2_6_port);
   y_i_6 : NAND2_28 port map( a => s1_6_port, b => s2_6_port, f => Y(6));
   s1_i_7 : NAND2_27 port map( a => A(7), b => sel_not, f => s1_7_port);
   s2_i_7 : NAND2_26 port map( a => B(7), b => SEL, f => s2_7_port);
   y_i_7 : NAND2_25 port map( a => s1_7_port, b => s2_7_port, f => Y(7));
   s1_i_8 : NAND2_24 port map( a => A(8), b => sel_not, f => s1_8_port);
   s2_i_8 : NAND2_23 port map( a => B(8), b => SEL, f => s2_8_port);
   y_i_8 : NAND2_22 port map( a => s1_8_port, b => s2_8_port, f => Y(8));
   s1_i_9 : NAND2_21 port map( a => A(9), b => sel_not, f => s1_9_port);
   s2_i_9 : NAND2_20 port map( a => B(9), b => SEL, f => s2_9_port);
   y_i_9 : NAND2_19 port map( a => s1_9_port, b => s2_9_port, f => Y(9));
   s1_i_10 : NAND2_18 port map( a => A(10), b => sel_not, f => s1_10_port);
   s2_i_10 : NAND2_17 port map( a => B(10), b => SEL, f => s2_10_port);
   y_i_10 : NAND2_16 port map( a => s1_10_port, b => s2_10_port, f => Y(10));
   s1_i_11 : NAND2_15 port map( a => A(11), b => sel_not, f => s1_11_port);
   s2_i_11 : NAND2_14 port map( a => B(11), b => SEL, f => s2_11_port);
   y_i_11 : NAND2_13 port map( a => s1_11_port, b => s2_11_port, f => Y(11));
   s1_i_12 : NAND2_12 port map( a => A(12), b => sel_not, f => s1_12_port);
   s2_i_12 : NAND2_11 port map( a => B(12), b => SEL, f => s2_12_port);
   y_i_12 : NAND2_10 port map( a => s1_12_port, b => s2_12_port, f => Y(12));
   s1_i_13 : NAND2_9 port map( a => A(13), b => sel_not, f => s1_13_port);
   s2_i_13 : NAND2_8 port map( a => B(13), b => SEL, f => s2_13_port);
   y_i_13 : NAND2_7 port map( a => s1_13_port, b => s2_13_port, f => Y(13));
   s1_i_14 : NAND2_6 port map( a => A(14), b => sel_not, f => s1_14_port);
   s2_i_14 : NAND2_5 port map( a => B(14), b => SEL, f => s2_14_port);
   y_i_14 : NAND2_4 port map( a => s1_14_port, b => s2_14_port, f => Y(14));
   s1_i_15 : NAND2_3 port map( a => A(15), b => sel_not, f => s1_15_port);
   s2_i_15 : NAND2_2 port map( a => B(15), b => SEL, f => s2_15_port);
   y_i_15 : NAND2_1 port map( a => s1_15_port, b => s2_15_port, f => Y(15));

end SYN_structural;
