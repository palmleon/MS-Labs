
library IEEE;

use IEEE.std_logic_1164.all;

package CONV_PACK_ACC_N64_1 is

-- define attributes
attribute ENUM_ENCODING : STRING;

end CONV_PACK_ACC_N64_1;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_63 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_63;

architecture SYN_ASYNCHARCH_EN of FD_63 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1000 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1000);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_62 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_62;

architecture SYN_ASYNCHARCH_EN of FD_62 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1001 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1001);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_61 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_61;

architecture SYN_ASYNCHARCH_EN of FD_61 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1002 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1002);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_60 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_60;

architecture SYN_ASYNCHARCH_EN of FD_60 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1003 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1003);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_59 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_59;

architecture SYN_ASYNCHARCH_EN of FD_59 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1004 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1004);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_58 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_58;

architecture SYN_ASYNCHARCH_EN of FD_58 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1005 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1005);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_57 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_57;

architecture SYN_ASYNCHARCH_EN of FD_57 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1006 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1006);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_56 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_56;

architecture SYN_ASYNCHARCH_EN of FD_56 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1007 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1007);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_55 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_55;

architecture SYN_ASYNCHARCH_EN of FD_55 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1008 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1008);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_54 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_54;

architecture SYN_ASYNCHARCH_EN of FD_54 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1009 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1009);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_53 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_53;

architecture SYN_ASYNCHARCH_EN of FD_53 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1010 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1010);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_52 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_52;

architecture SYN_ASYNCHARCH_EN of FD_52 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1011 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1011);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_51 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_51;

architecture SYN_ASYNCHARCH_EN of FD_51 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1012 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1012);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_50 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_50;

architecture SYN_ASYNCHARCH_EN of FD_50 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1013 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1013);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_49 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_49;

architecture SYN_ASYNCHARCH_EN of FD_49 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1014 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1014);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_48 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_48;

architecture SYN_ASYNCHARCH_EN of FD_48 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1015 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1015);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_47 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_47;

architecture SYN_ASYNCHARCH_EN of FD_47 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1016 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1016);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_46 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_46;

architecture SYN_ASYNCHARCH_EN of FD_46 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1017 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1017);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_45 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_45;

architecture SYN_ASYNCHARCH_EN of FD_45 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1018 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1018);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_44 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_44;

architecture SYN_ASYNCHARCH_EN of FD_44 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1019 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1019);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_43 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_43;

architecture SYN_ASYNCHARCH_EN of FD_43 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1020 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1020);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_42 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_42;

architecture SYN_ASYNCHARCH_EN of FD_42 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1021 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1021);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_41 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_41;

architecture SYN_ASYNCHARCH_EN of FD_41 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1022 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1022);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_40 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_40;

architecture SYN_ASYNCHARCH_EN of FD_40 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1023 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1023);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_39 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_39;

architecture SYN_ASYNCHARCH_EN of FD_39 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1024 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1024);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_38 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_38;

architecture SYN_ASYNCHARCH_EN of FD_38 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1025 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1025);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_37 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_37;

architecture SYN_ASYNCHARCH_EN of FD_37 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1026 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1026);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_36 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_36;

architecture SYN_ASYNCHARCH_EN of FD_36 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1027 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1027);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_35 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_35;

architecture SYN_ASYNCHARCH_EN of FD_35 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1028 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1028);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_34 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_34;

architecture SYN_ASYNCHARCH_EN of FD_34 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1029 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1029);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_33 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_33;

architecture SYN_ASYNCHARCH_EN of FD_33 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1030 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1030);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_32 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_32;

architecture SYN_ASYNCHARCH_EN of FD_32 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1031 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1031);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_31 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_31;

architecture SYN_ASYNCHARCH_EN of FD_31 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1032 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1032);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_30 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_30;

architecture SYN_ASYNCHARCH_EN of FD_30 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1033 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1033);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_29 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_29;

architecture SYN_ASYNCHARCH_EN of FD_29 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1034 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1034);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_28 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_28;

architecture SYN_ASYNCHARCH_EN of FD_28 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1035 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1035);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_27 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_27;

architecture SYN_ASYNCHARCH_EN of FD_27 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1036 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1036);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_26 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_26;

architecture SYN_ASYNCHARCH_EN of FD_26 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1037 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1037);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_25 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_25;

architecture SYN_ASYNCHARCH_EN of FD_25 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1038 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1038);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_24 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_24;

architecture SYN_ASYNCHARCH_EN of FD_24 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1039 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1039);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_23 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_23;

architecture SYN_ASYNCHARCH_EN of FD_23 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1040 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1040);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_22 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_22;

architecture SYN_ASYNCHARCH_EN of FD_22 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1041 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1041);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_21 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_21;

architecture SYN_ASYNCHARCH_EN of FD_21 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1042 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1042);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_20 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_20;

architecture SYN_ASYNCHARCH_EN of FD_20 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1043 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1043);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_19 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_19;

architecture SYN_ASYNCHARCH_EN of FD_19 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1044 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1044);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_18 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_18;

architecture SYN_ASYNCHARCH_EN of FD_18 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1045 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1045);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_17 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_17;

architecture SYN_ASYNCHARCH_EN of FD_17 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1046 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1046);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_16 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_16;

architecture SYN_ASYNCHARCH_EN of FD_16 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1047 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1047);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_15 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_15;

architecture SYN_ASYNCHARCH_EN of FD_15 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1048 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1048);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_14 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_14;

architecture SYN_ASYNCHARCH_EN of FD_14 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1049 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1049);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_13 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_13;

architecture SYN_ASYNCHARCH_EN of FD_13 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1050 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1050);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_12 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_12;

architecture SYN_ASYNCHARCH_EN of FD_12 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1051 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1051);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_11 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_11;

architecture SYN_ASYNCHARCH_EN of FD_11 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1052 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1052);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_10 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_10;

architecture SYN_ASYNCHARCH_EN of FD_10 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1053 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1053);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_9 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_9;

architecture SYN_ASYNCHARCH_EN of FD_9 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1054 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1054);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_8 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_8;

architecture SYN_ASYNCHARCH_EN of FD_8 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1055 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1055);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_7 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_7;

architecture SYN_ASYNCHARCH_EN of FD_7 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1056 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1056);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_6 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_6;

architecture SYN_ASYNCHARCH_EN of FD_6 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1057 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1057);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_5 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_5;

architecture SYN_ASYNCHARCH_EN of FD_5 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1058 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1058);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_4 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_4;

architecture SYN_ASYNCHARCH_EN of FD_4 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1059 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1059);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_3 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_3;

architecture SYN_ASYNCHARCH_EN of FD_3 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1060 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1060);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_2 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_2;

architecture SYN_ASYNCHARCH_EN of FD_2 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1061 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1061);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_1 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_1;

architecture SYN_ASYNCHARCH_EN of FD_1 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n1, n2, n_1062 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n1, CK => CK, RN => n2, Q => Q_port, QN => 
                           n_1062);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n1);
   U3 : INV_X1 port map( A => RESET, ZN => n2);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_63 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_63;

architecture SYN_BEHAVIORAL of FA_63 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_62 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_62;

architecture SYN_BEHAVIORAL of FA_62 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_61 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_61;

architecture SYN_BEHAVIORAL of FA_61 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_60 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_60;

architecture SYN_BEHAVIORAL of FA_60 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_59 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_59;

architecture SYN_BEHAVIORAL of FA_59 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_58 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_58;

architecture SYN_BEHAVIORAL of FA_58 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_57 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_57;

architecture SYN_BEHAVIORAL of FA_57 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_56 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_56;

architecture SYN_BEHAVIORAL of FA_56 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_55 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_55;

architecture SYN_BEHAVIORAL of FA_55 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_54 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_54;

architecture SYN_BEHAVIORAL of FA_54 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_53 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_53;

architecture SYN_BEHAVIORAL of FA_53 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_52 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_52;

architecture SYN_BEHAVIORAL of FA_52 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_51 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_51;

architecture SYN_BEHAVIORAL of FA_51 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_50 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_50;

architecture SYN_BEHAVIORAL of FA_50 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_49 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_49;

architecture SYN_BEHAVIORAL of FA_49 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_48 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_48;

architecture SYN_BEHAVIORAL of FA_48 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_47 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_47;

architecture SYN_BEHAVIORAL of FA_47 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_46 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_46;

architecture SYN_BEHAVIORAL of FA_46 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_45 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_45;

architecture SYN_BEHAVIORAL of FA_45 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_44 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_44;

architecture SYN_BEHAVIORAL of FA_44 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_43 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_43;

architecture SYN_BEHAVIORAL of FA_43 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_42 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_42;

architecture SYN_BEHAVIORAL of FA_42 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_41 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_41;

architecture SYN_BEHAVIORAL of FA_41 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_40 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_40;

architecture SYN_BEHAVIORAL of FA_40 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_39 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_39;

architecture SYN_BEHAVIORAL of FA_39 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_38 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_38;

architecture SYN_BEHAVIORAL of FA_38 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_37 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_37;

architecture SYN_BEHAVIORAL of FA_37 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_36 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_36;

architecture SYN_BEHAVIORAL of FA_36 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_35 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_35;

architecture SYN_BEHAVIORAL of FA_35 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_34 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_34;

architecture SYN_BEHAVIORAL of FA_34 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_33 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_33;

architecture SYN_BEHAVIORAL of FA_33 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_32 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_32;

architecture SYN_BEHAVIORAL of FA_32 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_31 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_31;

architecture SYN_BEHAVIORAL of FA_31 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_30 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_30;

architecture SYN_BEHAVIORAL of FA_30 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_29 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_29;

architecture SYN_BEHAVIORAL of FA_29 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_28 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_28;

architecture SYN_BEHAVIORAL of FA_28 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_27 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_27;

architecture SYN_BEHAVIORAL of FA_27 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_26 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_26;

architecture SYN_BEHAVIORAL of FA_26 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_25 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_25;

architecture SYN_BEHAVIORAL of FA_25 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_24 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_24;

architecture SYN_BEHAVIORAL of FA_24 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_23 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_23;

architecture SYN_BEHAVIORAL of FA_23 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_22 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_22;

architecture SYN_BEHAVIORAL of FA_22 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_21 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_21;

architecture SYN_BEHAVIORAL of FA_21 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_20 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_20;

architecture SYN_BEHAVIORAL of FA_20 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_19 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_19;

architecture SYN_BEHAVIORAL of FA_19 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_18 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_18;

architecture SYN_BEHAVIORAL of FA_18 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_17 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_17;

architecture SYN_BEHAVIORAL of FA_17 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_16 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_16;

architecture SYN_BEHAVIORAL of FA_16 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_15 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_15;

architecture SYN_BEHAVIORAL of FA_15 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_14 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_14;

architecture SYN_BEHAVIORAL of FA_14 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_13 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_13;

architecture SYN_BEHAVIORAL of FA_13 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_12 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_12;

architecture SYN_BEHAVIORAL of FA_12 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_11 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_11;

architecture SYN_BEHAVIORAL of FA_11 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_10 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_10;

architecture SYN_BEHAVIORAL of FA_10 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_9 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_9;

architecture SYN_BEHAVIORAL of FA_9 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_8 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_8;

architecture SYN_BEHAVIORAL of FA_8 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_7 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_7;

architecture SYN_BEHAVIORAL of FA_7 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_6 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_6;

architecture SYN_BEHAVIORAL of FA_6 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_5 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_5;

architecture SYN_BEHAVIORAL of FA_5 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_4 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_4;

architecture SYN_BEHAVIORAL of FA_4 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_3 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_3;

architecture SYN_BEHAVIORAL of FA_3 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_2 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_2;

architecture SYN_BEHAVIORAL of FA_2 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_1 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_1;

architecture SYN_BEHAVIORAL of FA_1 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_191 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_191;

architecture SYN_behavioral of NAND2_191 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_190 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_190;

architecture SYN_behavioral of NAND2_190 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_189 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_189;

architecture SYN_behavioral of NAND2_189 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_188 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_188;

architecture SYN_behavioral of NAND2_188 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_187 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_187;

architecture SYN_behavioral of NAND2_187 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_186 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_186;

architecture SYN_behavioral of NAND2_186 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_185 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_185;

architecture SYN_behavioral of NAND2_185 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_184 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_184;

architecture SYN_behavioral of NAND2_184 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_183 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_183;

architecture SYN_behavioral of NAND2_183 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_182 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_182;

architecture SYN_behavioral of NAND2_182 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_181 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_181;

architecture SYN_behavioral of NAND2_181 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_180 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_180;

architecture SYN_behavioral of NAND2_180 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_179 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_179;

architecture SYN_behavioral of NAND2_179 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_178 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_178;

architecture SYN_behavioral of NAND2_178 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_177 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_177;

architecture SYN_behavioral of NAND2_177 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_176 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_176;

architecture SYN_behavioral of NAND2_176 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_175 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_175;

architecture SYN_behavioral of NAND2_175 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_174 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_174;

architecture SYN_behavioral of NAND2_174 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_173 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_173;

architecture SYN_behavioral of NAND2_173 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_172 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_172;

architecture SYN_behavioral of NAND2_172 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_171 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_171;

architecture SYN_behavioral of NAND2_171 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_170 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_170;

architecture SYN_behavioral of NAND2_170 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_169 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_169;

architecture SYN_behavioral of NAND2_169 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_168 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_168;

architecture SYN_behavioral of NAND2_168 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_167 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_167;

architecture SYN_behavioral of NAND2_167 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_166 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_166;

architecture SYN_behavioral of NAND2_166 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_165 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_165;

architecture SYN_behavioral of NAND2_165 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_164 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_164;

architecture SYN_behavioral of NAND2_164 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_163 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_163;

architecture SYN_behavioral of NAND2_163 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_162 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_162;

architecture SYN_behavioral of NAND2_162 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_161 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_161;

architecture SYN_behavioral of NAND2_161 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_160 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_160;

architecture SYN_behavioral of NAND2_160 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_159 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_159;

architecture SYN_behavioral of NAND2_159 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_158 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_158;

architecture SYN_behavioral of NAND2_158 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_157 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_157;

architecture SYN_behavioral of NAND2_157 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_156 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_156;

architecture SYN_behavioral of NAND2_156 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_155 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_155;

architecture SYN_behavioral of NAND2_155 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_154 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_154;

architecture SYN_behavioral of NAND2_154 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_153 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_153;

architecture SYN_behavioral of NAND2_153 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_152 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_152;

architecture SYN_behavioral of NAND2_152 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_151 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_151;

architecture SYN_behavioral of NAND2_151 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_150 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_150;

architecture SYN_behavioral of NAND2_150 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_149 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_149;

architecture SYN_behavioral of NAND2_149 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_148 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_148;

architecture SYN_behavioral of NAND2_148 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_147 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_147;

architecture SYN_behavioral of NAND2_147 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_146 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_146;

architecture SYN_behavioral of NAND2_146 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_145 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_145;

architecture SYN_behavioral of NAND2_145 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_144 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_144;

architecture SYN_behavioral of NAND2_144 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_143 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_143;

architecture SYN_behavioral of NAND2_143 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_142 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_142;

architecture SYN_behavioral of NAND2_142 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_141 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_141;

architecture SYN_behavioral of NAND2_141 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_140 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_140;

architecture SYN_behavioral of NAND2_140 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_139 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_139;

architecture SYN_behavioral of NAND2_139 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_138 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_138;

architecture SYN_behavioral of NAND2_138 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_137 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_137;

architecture SYN_behavioral of NAND2_137 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_136 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_136;

architecture SYN_behavioral of NAND2_136 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_135 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_135;

architecture SYN_behavioral of NAND2_135 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_134 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_134;

architecture SYN_behavioral of NAND2_134 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_133 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_133;

architecture SYN_behavioral of NAND2_133 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_132 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_132;

architecture SYN_behavioral of NAND2_132 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_131 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_131;

architecture SYN_behavioral of NAND2_131 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_130 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_130;

architecture SYN_behavioral of NAND2_130 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_129 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_129;

architecture SYN_behavioral of NAND2_129 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_128 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_128;

architecture SYN_behavioral of NAND2_128 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_127 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_127;

architecture SYN_behavioral of NAND2_127 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_126 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_126;

architecture SYN_behavioral of NAND2_126 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_125 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_125;

architecture SYN_behavioral of NAND2_125 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_124 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_124;

architecture SYN_behavioral of NAND2_124 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_123 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_123;

architecture SYN_behavioral of NAND2_123 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_122 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_122;

architecture SYN_behavioral of NAND2_122 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_121 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_121;

architecture SYN_behavioral of NAND2_121 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_120 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_120;

architecture SYN_behavioral of NAND2_120 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_119 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_119;

architecture SYN_behavioral of NAND2_119 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_118 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_118;

architecture SYN_behavioral of NAND2_118 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_117 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_117;

architecture SYN_behavioral of NAND2_117 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_116 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_116;

architecture SYN_behavioral of NAND2_116 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_115 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_115;

architecture SYN_behavioral of NAND2_115 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_114 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_114;

architecture SYN_behavioral of NAND2_114 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_113 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_113;

architecture SYN_behavioral of NAND2_113 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_112 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_112;

architecture SYN_behavioral of NAND2_112 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_111 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_111;

architecture SYN_behavioral of NAND2_111 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_110 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_110;

architecture SYN_behavioral of NAND2_110 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_109 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_109;

architecture SYN_behavioral of NAND2_109 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_108 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_108;

architecture SYN_behavioral of NAND2_108 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_107 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_107;

architecture SYN_behavioral of NAND2_107 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_106 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_106;

architecture SYN_behavioral of NAND2_106 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_105 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_105;

architecture SYN_behavioral of NAND2_105 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_104 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_104;

architecture SYN_behavioral of NAND2_104 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_103 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_103;

architecture SYN_behavioral of NAND2_103 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_102 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_102;

architecture SYN_behavioral of NAND2_102 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_101 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_101;

architecture SYN_behavioral of NAND2_101 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_100 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_100;

architecture SYN_behavioral of NAND2_100 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_99 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_99;

architecture SYN_behavioral of NAND2_99 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_98 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_98;

architecture SYN_behavioral of NAND2_98 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_97 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_97;

architecture SYN_behavioral of NAND2_97 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_96 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_96;

architecture SYN_behavioral of NAND2_96 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_95 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_95;

architecture SYN_behavioral of NAND2_95 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_94 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_94;

architecture SYN_behavioral of NAND2_94 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_93 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_93;

architecture SYN_behavioral of NAND2_93 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_92 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_92;

architecture SYN_behavioral of NAND2_92 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_91 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_91;

architecture SYN_behavioral of NAND2_91 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_90 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_90;

architecture SYN_behavioral of NAND2_90 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_89 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_89;

architecture SYN_behavioral of NAND2_89 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_88 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_88;

architecture SYN_behavioral of NAND2_88 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_87 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_87;

architecture SYN_behavioral of NAND2_87 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_86 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_86;

architecture SYN_behavioral of NAND2_86 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_85 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_85;

architecture SYN_behavioral of NAND2_85 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_84 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_84;

architecture SYN_behavioral of NAND2_84 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_83 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_83;

architecture SYN_behavioral of NAND2_83 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_82 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_82;

architecture SYN_behavioral of NAND2_82 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_81 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_81;

architecture SYN_behavioral of NAND2_81 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_80 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_80;

architecture SYN_behavioral of NAND2_80 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_79 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_79;

architecture SYN_behavioral of NAND2_79 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_78 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_78;

architecture SYN_behavioral of NAND2_78 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_77 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_77;

architecture SYN_behavioral of NAND2_77 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_76 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_76;

architecture SYN_behavioral of NAND2_76 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_75 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_75;

architecture SYN_behavioral of NAND2_75 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_74 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_74;

architecture SYN_behavioral of NAND2_74 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_73 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_73;

architecture SYN_behavioral of NAND2_73 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_72 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_72;

architecture SYN_behavioral of NAND2_72 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_71 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_71;

architecture SYN_behavioral of NAND2_71 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_70 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_70;

architecture SYN_behavioral of NAND2_70 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_69 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_69;

architecture SYN_behavioral of NAND2_69 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_68 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_68;

architecture SYN_behavioral of NAND2_68 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_67 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_67;

architecture SYN_behavioral of NAND2_67 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_66 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_66;

architecture SYN_behavioral of NAND2_66 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_65 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_65;

architecture SYN_behavioral of NAND2_65 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_64 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_64;

architecture SYN_behavioral of NAND2_64 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_63 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_63;

architecture SYN_behavioral of NAND2_63 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_62 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_62;

architecture SYN_behavioral of NAND2_62 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_61 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_61;

architecture SYN_behavioral of NAND2_61 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_60 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_60;

architecture SYN_behavioral of NAND2_60 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_59 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_59;

architecture SYN_behavioral of NAND2_59 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_58 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_58;

architecture SYN_behavioral of NAND2_58 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_57 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_57;

architecture SYN_behavioral of NAND2_57 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_56 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_56;

architecture SYN_behavioral of NAND2_56 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_55 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_55;

architecture SYN_behavioral of NAND2_55 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_54 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_54;

architecture SYN_behavioral of NAND2_54 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_53 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_53;

architecture SYN_behavioral of NAND2_53 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_52 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_52;

architecture SYN_behavioral of NAND2_52 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_51 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_51;

architecture SYN_behavioral of NAND2_51 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_50 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_50;

architecture SYN_behavioral of NAND2_50 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_49 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_49;

architecture SYN_behavioral of NAND2_49 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_48 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_48;

architecture SYN_behavioral of NAND2_48 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_47 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_47;

architecture SYN_behavioral of NAND2_47 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_46 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_46;

architecture SYN_behavioral of NAND2_46 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_45 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_45;

architecture SYN_behavioral of NAND2_45 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_44 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_44;

architecture SYN_behavioral of NAND2_44 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_43 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_43;

architecture SYN_behavioral of NAND2_43 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_42 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_42;

architecture SYN_behavioral of NAND2_42 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_41 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_41;

architecture SYN_behavioral of NAND2_41 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_40 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_40;

architecture SYN_behavioral of NAND2_40 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_39 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_39;

architecture SYN_behavioral of NAND2_39 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_38 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_38;

architecture SYN_behavioral of NAND2_38 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_37 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_37;

architecture SYN_behavioral of NAND2_37 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_36 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_36;

architecture SYN_behavioral of NAND2_36 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_35 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_35;

architecture SYN_behavioral of NAND2_35 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_34 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_34;

architecture SYN_behavioral of NAND2_34 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_33 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_33;

architecture SYN_behavioral of NAND2_33 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_32 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_32;

architecture SYN_behavioral of NAND2_32 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_31 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_31;

architecture SYN_behavioral of NAND2_31 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_30 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_30;

architecture SYN_behavioral of NAND2_30 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_29 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_29;

architecture SYN_behavioral of NAND2_29 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_28 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_28;

architecture SYN_behavioral of NAND2_28 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_27 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_27;

architecture SYN_behavioral of NAND2_27 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_26 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_26;

architecture SYN_behavioral of NAND2_26 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_25 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_25;

architecture SYN_behavioral of NAND2_25 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_24 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_24;

architecture SYN_behavioral of NAND2_24 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_23 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_23;

architecture SYN_behavioral of NAND2_23 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_22 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_22;

architecture SYN_behavioral of NAND2_22 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_21 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_21;

architecture SYN_behavioral of NAND2_21 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_20 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_20;

architecture SYN_behavioral of NAND2_20 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_19 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_19;

architecture SYN_behavioral of NAND2_19 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_18 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_18;

architecture SYN_behavioral of NAND2_18 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_17 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_17;

architecture SYN_behavioral of NAND2_17 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_16 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_16;

architecture SYN_behavioral of NAND2_16 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_15 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_15;

architecture SYN_behavioral of NAND2_15 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_14 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_14;

architecture SYN_behavioral of NAND2_14 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_13 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_13;

architecture SYN_behavioral of NAND2_13 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_12 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_12;

architecture SYN_behavioral of NAND2_12 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_11 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_11;

architecture SYN_behavioral of NAND2_11 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_10 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_10;

architecture SYN_behavioral of NAND2_10 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_9 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_9;

architecture SYN_behavioral of NAND2_9 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_8 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_8;

architecture SYN_behavioral of NAND2_8 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_7 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_7;

architecture SYN_behavioral of NAND2_7 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_6 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_6;

architecture SYN_behavioral of NAND2_6 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_5 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_5;

architecture SYN_behavioral of NAND2_5 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_4 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_4;

architecture SYN_behavioral of NAND2_4 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_3 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_3;

architecture SYN_behavioral of NAND2_3 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_2 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_2;

architecture SYN_behavioral of NAND2_2 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_1 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_1;

architecture SYN_behavioral of NAND2_1 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_0 is

   port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);

end FD_0;

architecture SYN_ASYNCHARCH_EN of FD_0 is

   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component MUX2_X1
      port( A, B, S : in std_logic;  Z : out std_logic);
   end component;
   
   component DFFR_X1
      port( D, CK, RN : in std_logic;  Q, QN : out std_logic);
   end component;
   
   signal Q_port, n3, n4, n_1063 : std_logic;

begin
   Q <= Q_port;
   
   Q_reg : DFFR_X1 port map( D => n4, CK => CK, RN => n3, Q => Q_port, QN => 
                           n_1063);
   U2 : MUX2_X1 port map( A => Q_port, B => D, S => ENABLE, Z => n4);
   U3 : INV_X1 port map( A => RESET, ZN => n3);

end SYN_ASYNCHARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FA_0 is

   port( A, B, Ci : in std_logic;  S, Co : out std_logic);

end FA_0;

architecture SYN_BEHAVIORAL of FA_0 is

   component XOR2_X1
      port( A, B : in std_logic;  Z : out std_logic);
   end component;
   
   component AOI22_X1
      port( A1, A2, B1, B2 : in std_logic;  ZN : out std_logic);
   end component;
   
   component INV_X1
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   signal n1, n2 : std_logic;

begin
   
   U1 : XOR2_X1 port map( A => Ci, B => n1, Z => S);
   U2 : INV_X1 port map( A => n2, ZN => Co);
   U3 : AOI22_X1 port map( A1 => B, A2 => A, B1 => n1, B2 => Ci, ZN => n2);
   U4 : XOR2_X1 port map( A => A, B => B, Z => n1);

end SYN_BEHAVIORAL;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity NAND2_0 is

   port( a, b : in std_logic;  f : out std_logic);

end NAND2_0;

architecture SYN_behavioral of NAND2_0 is

   component NAND2_X1
      port( A1, A2 : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : NAND2_X1 port map( A1 => b, A2 => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity INV is

   port( a : in std_logic;  f : out std_logic);

end INV;

architecture SYN_behavioral of INV is

   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;

begin
   
   U1 : INV_X4 port map( A => a, ZN => f);

end SYN_behavioral;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity FD_GENERIC_N64 is

   port( D : in std_logic_vector (63 downto 0);  CK, RESET, ENABLE : in 
         std_logic;  Q : out std_logic_vector (63 downto 0));

end FD_GENERIC_N64;

architecture SYN_ASYNCARCH_EN of FD_GENERIC_N64 is

   component FD_1
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_2
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_3
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_4
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_5
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_6
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_7
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_8
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_9
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_10
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_11
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_12
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_13
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_14
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_15
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_16
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_17
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_18
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_19
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_20
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_21
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_22
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_23
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_24
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_25
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_26
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_27
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_28
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_29
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_30
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_31
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_32
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_33
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_34
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_35
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_36
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_37
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_38
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_39
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_40
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_41
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_42
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_43
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_44
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_45
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_46
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_47
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_48
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_49
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_50
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_51
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_52
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_53
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_54
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_55
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_56
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_57
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_58
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_59
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_60
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_61
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_62
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_63
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;
   
   component FD_0
      port( D, CK, RESET, ENABLE : in std_logic;  Q : out std_logic);
   end component;

begin
   
   FF_0 : FD_0 port map( D => D(0), CK => CK, RESET => RESET, ENABLE => ENABLE,
                           Q => Q(0));
   FF_1 : FD_63 port map( D => D(1), CK => CK, RESET => RESET, ENABLE => ENABLE
                           , Q => Q(1));
   FF_2 : FD_62 port map( D => D(2), CK => CK, RESET => RESET, ENABLE => ENABLE
                           , Q => Q(2));
   FF_3 : FD_61 port map( D => D(3), CK => CK, RESET => RESET, ENABLE => ENABLE
                           , Q => Q(3));
   FF_4 : FD_60 port map( D => D(4), CK => CK, RESET => RESET, ENABLE => ENABLE
                           , Q => Q(4));
   FF_5 : FD_59 port map( D => D(5), CK => CK, RESET => RESET, ENABLE => ENABLE
                           , Q => Q(5));
   FF_6 : FD_58 port map( D => D(6), CK => CK, RESET => RESET, ENABLE => ENABLE
                           , Q => Q(6));
   FF_7 : FD_57 port map( D => D(7), CK => CK, RESET => RESET, ENABLE => ENABLE
                           , Q => Q(7));
   FF_8 : FD_56 port map( D => D(8), CK => CK, RESET => RESET, ENABLE => ENABLE
                           , Q => Q(8));
   FF_9 : FD_55 port map( D => D(9), CK => CK, RESET => RESET, ENABLE => ENABLE
                           , Q => Q(9));
   FF_10 : FD_54 port map( D => D(10), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(10));
   FF_11 : FD_53 port map( D => D(11), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(11));
   FF_12 : FD_52 port map( D => D(12), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(12));
   FF_13 : FD_51 port map( D => D(13), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(13));
   FF_14 : FD_50 port map( D => D(14), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(14));
   FF_15 : FD_49 port map( D => D(15), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(15));
   FF_16 : FD_48 port map( D => D(16), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(16));
   FF_17 : FD_47 port map( D => D(17), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(17));
   FF_18 : FD_46 port map( D => D(18), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(18));
   FF_19 : FD_45 port map( D => D(19), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(19));
   FF_20 : FD_44 port map( D => D(20), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(20));
   FF_21 : FD_43 port map( D => D(21), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(21));
   FF_22 : FD_42 port map( D => D(22), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(22));
   FF_23 : FD_41 port map( D => D(23), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(23));
   FF_24 : FD_40 port map( D => D(24), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(24));
   FF_25 : FD_39 port map( D => D(25), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(25));
   FF_26 : FD_38 port map( D => D(26), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(26));
   FF_27 : FD_37 port map( D => D(27), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(27));
   FF_28 : FD_36 port map( D => D(28), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(28));
   FF_29 : FD_35 port map( D => D(29), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(29));
   FF_30 : FD_34 port map( D => D(30), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(30));
   FF_31 : FD_33 port map( D => D(31), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(31));
   FF_32 : FD_32 port map( D => D(32), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(32));
   FF_33 : FD_31 port map( D => D(33), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(33));
   FF_34 : FD_30 port map( D => D(34), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(34));
   FF_35 : FD_29 port map( D => D(35), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(35));
   FF_36 : FD_28 port map( D => D(36), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(36));
   FF_37 : FD_27 port map( D => D(37), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(37));
   FF_38 : FD_26 port map( D => D(38), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(38));
   FF_39 : FD_25 port map( D => D(39), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(39));
   FF_40 : FD_24 port map( D => D(40), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(40));
   FF_41 : FD_23 port map( D => D(41), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(41));
   FF_42 : FD_22 port map( D => D(42), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(42));
   FF_43 : FD_21 port map( D => D(43), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(43));
   FF_44 : FD_20 port map( D => D(44), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(44));
   FF_45 : FD_19 port map( D => D(45), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(45));
   FF_46 : FD_18 port map( D => D(46), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(46));
   FF_47 : FD_17 port map( D => D(47), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(47));
   FF_48 : FD_16 port map( D => D(48), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(48));
   FF_49 : FD_15 port map( D => D(49), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(49));
   FF_50 : FD_14 port map( D => D(50), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(50));
   FF_51 : FD_13 port map( D => D(51), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(51));
   FF_52 : FD_12 port map( D => D(52), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(52));
   FF_53 : FD_11 port map( D => D(53), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(53));
   FF_54 : FD_10 port map( D => D(54), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(54));
   FF_55 : FD_9 port map( D => D(55), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(55));
   FF_56 : FD_8 port map( D => D(56), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(56));
   FF_57 : FD_7 port map( D => D(57), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(57));
   FF_58 : FD_6 port map( D => D(58), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(58));
   FF_59 : FD_5 port map( D => D(59), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(59));
   FF_60 : FD_4 port map( D => D(60), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(60));
   FF_61 : FD_3 port map( D => D(61), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(61));
   FF_62 : FD_2 port map( D => D(62), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(62));
   FF_63 : FD_1 port map( D => D(63), CK => CK, RESET => RESET, ENABLE => 
                           ENABLE, Q => Q(63));

end SYN_ASYNCARCH_EN;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity RCA_N64 is

   port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : out
         std_logic_vector (63 downto 0);  Co : out std_logic);

end RCA_N64;

architecture SYN_structural of RCA_N64 is

   component FA_1
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_2
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_3
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_4
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_5
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_6
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_7
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_8
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_9
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_10
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_11
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_12
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_13
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_14
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_15
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_16
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_17
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_18
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_19
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_20
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_21
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_22
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_23
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_24
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_25
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_26
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_27
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_28
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_29
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_30
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_31
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_32
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_33
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_34
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_35
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_36
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_37
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_38
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_39
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_40
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_41
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_42
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_43
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_44
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_45
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_46
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_47
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_48
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_49
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_50
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_51
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_52
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_53
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_54
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_55
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_56
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_57
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_58
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_59
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_60
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_61
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_62
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_63
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   component FA_0
      port( A, B, Ci : in std_logic;  S, Co : out std_logic);
   end component;
   
   signal tmp_63_port, tmp_62_port, tmp_61_port, tmp_60_port, tmp_59_port, 
      tmp_58_port, tmp_57_port, tmp_56_port, tmp_55_port, tmp_54_port, 
      tmp_53_port, tmp_52_port, tmp_51_port, tmp_50_port, tmp_49_port, 
      tmp_48_port, tmp_47_port, tmp_46_port, tmp_45_port, tmp_44_port, 
      tmp_43_port, tmp_42_port, tmp_41_port, tmp_40_port, tmp_39_port, 
      tmp_38_port, tmp_37_port, tmp_36_port, tmp_35_port, tmp_34_port, 
      tmp_33_port, tmp_32_port, tmp_31_port, tmp_30_port, tmp_29_port, 
      tmp_28_port, tmp_27_port, tmp_26_port, tmp_25_port, tmp_24_port, 
      tmp_23_port, tmp_22_port, tmp_21_port, tmp_20_port, tmp_19_port, 
      tmp_18_port, tmp_17_port, tmp_16_port, tmp_15_port, tmp_14_port, 
      tmp_13_port, tmp_12_port, tmp_11_port, tmp_10_port, tmp_9_port, 
      tmp_8_port, tmp_7_port, tmp_6_port, tmp_5_port, tmp_4_port, tmp_3_port, 
      tmp_2_port, tmp_1_port : std_logic;

begin
   
   FAi_0 : FA_0 port map( A => A(0), B => B(0), Ci => Ci, S => S(0), Co => 
                           tmp_1_port);
   FAi_1 : FA_63 port map( A => A(1), B => B(1), Ci => tmp_1_port, S => S(1), 
                           Co => tmp_2_port);
   FAi_2 : FA_62 port map( A => A(2), B => B(2), Ci => tmp_2_port, S => S(2), 
                           Co => tmp_3_port);
   FAi_3 : FA_61 port map( A => A(3), B => B(3), Ci => tmp_3_port, S => S(3), 
                           Co => tmp_4_port);
   FAi_4 : FA_60 port map( A => A(4), B => B(4), Ci => tmp_4_port, S => S(4), 
                           Co => tmp_5_port);
   FAi_5 : FA_59 port map( A => A(5), B => B(5), Ci => tmp_5_port, S => S(5), 
                           Co => tmp_6_port);
   FAi_6 : FA_58 port map( A => A(6), B => B(6), Ci => tmp_6_port, S => S(6), 
                           Co => tmp_7_port);
   FAi_7 : FA_57 port map( A => A(7), B => B(7), Ci => tmp_7_port, S => S(7), 
                           Co => tmp_8_port);
   FAi_8 : FA_56 port map( A => A(8), B => B(8), Ci => tmp_8_port, S => S(8), 
                           Co => tmp_9_port);
   FAi_9 : FA_55 port map( A => A(9), B => B(9), Ci => tmp_9_port, S => S(9), 
                           Co => tmp_10_port);
   FAi_10 : FA_54 port map( A => A(10), B => B(10), Ci => tmp_10_port, S => 
                           S(10), Co => tmp_11_port);
   FAi_11 : FA_53 port map( A => A(11), B => B(11), Ci => tmp_11_port, S => 
                           S(11), Co => tmp_12_port);
   FAi_12 : FA_52 port map( A => A(12), B => B(12), Ci => tmp_12_port, S => 
                           S(12), Co => tmp_13_port);
   FAi_13 : FA_51 port map( A => A(13), B => B(13), Ci => tmp_13_port, S => 
                           S(13), Co => tmp_14_port);
   FAi_14 : FA_50 port map( A => A(14), B => B(14), Ci => tmp_14_port, S => 
                           S(14), Co => tmp_15_port);
   FAi_15 : FA_49 port map( A => A(15), B => B(15), Ci => tmp_15_port, S => 
                           S(15), Co => tmp_16_port);
   FAi_16 : FA_48 port map( A => A(16), B => B(16), Ci => tmp_16_port, S => 
                           S(16), Co => tmp_17_port);
   FAi_17 : FA_47 port map( A => A(17), B => B(17), Ci => tmp_17_port, S => 
                           S(17), Co => tmp_18_port);
   FAi_18 : FA_46 port map( A => A(18), B => B(18), Ci => tmp_18_port, S => 
                           S(18), Co => tmp_19_port);
   FAi_19 : FA_45 port map( A => A(19), B => B(19), Ci => tmp_19_port, S => 
                           S(19), Co => tmp_20_port);
   FAi_20 : FA_44 port map( A => A(20), B => B(20), Ci => tmp_20_port, S => 
                           S(20), Co => tmp_21_port);
   FAi_21 : FA_43 port map( A => A(21), B => B(21), Ci => tmp_21_port, S => 
                           S(21), Co => tmp_22_port);
   FAi_22 : FA_42 port map( A => A(22), B => B(22), Ci => tmp_22_port, S => 
                           S(22), Co => tmp_23_port);
   FAi_23 : FA_41 port map( A => A(23), B => B(23), Ci => tmp_23_port, S => 
                           S(23), Co => tmp_24_port);
   FAi_24 : FA_40 port map( A => A(24), B => B(24), Ci => tmp_24_port, S => 
                           S(24), Co => tmp_25_port);
   FAi_25 : FA_39 port map( A => A(25), B => B(25), Ci => tmp_25_port, S => 
                           S(25), Co => tmp_26_port);
   FAi_26 : FA_38 port map( A => A(26), B => B(26), Ci => tmp_26_port, S => 
                           S(26), Co => tmp_27_port);
   FAi_27 : FA_37 port map( A => A(27), B => B(27), Ci => tmp_27_port, S => 
                           S(27), Co => tmp_28_port);
   FAi_28 : FA_36 port map( A => A(28), B => B(28), Ci => tmp_28_port, S => 
                           S(28), Co => tmp_29_port);
   FAi_29 : FA_35 port map( A => A(29), B => B(29), Ci => tmp_29_port, S => 
                           S(29), Co => tmp_30_port);
   FAi_30 : FA_34 port map( A => A(30), B => B(30), Ci => tmp_30_port, S => 
                           S(30), Co => tmp_31_port);
   FAi_31 : FA_33 port map( A => A(31), B => B(31), Ci => tmp_31_port, S => 
                           S(31), Co => tmp_32_port);
   FAi_32 : FA_32 port map( A => A(32), B => B(32), Ci => tmp_32_port, S => 
                           S(32), Co => tmp_33_port);
   FAi_33 : FA_31 port map( A => A(33), B => B(33), Ci => tmp_33_port, S => 
                           S(33), Co => tmp_34_port);
   FAi_34 : FA_30 port map( A => A(34), B => B(34), Ci => tmp_34_port, S => 
                           S(34), Co => tmp_35_port);
   FAi_35 : FA_29 port map( A => A(35), B => B(35), Ci => tmp_35_port, S => 
                           S(35), Co => tmp_36_port);
   FAi_36 : FA_28 port map( A => A(36), B => B(36), Ci => tmp_36_port, S => 
                           S(36), Co => tmp_37_port);
   FAi_37 : FA_27 port map( A => A(37), B => B(37), Ci => tmp_37_port, S => 
                           S(37), Co => tmp_38_port);
   FAi_38 : FA_26 port map( A => A(38), B => B(38), Ci => tmp_38_port, S => 
                           S(38), Co => tmp_39_port);
   FAi_39 : FA_25 port map( A => A(39), B => B(39), Ci => tmp_39_port, S => 
                           S(39), Co => tmp_40_port);
   FAi_40 : FA_24 port map( A => A(40), B => B(40), Ci => tmp_40_port, S => 
                           S(40), Co => tmp_41_port);
   FAi_41 : FA_23 port map( A => A(41), B => B(41), Ci => tmp_41_port, S => 
                           S(41), Co => tmp_42_port);
   FAi_42 : FA_22 port map( A => A(42), B => B(42), Ci => tmp_42_port, S => 
                           S(42), Co => tmp_43_port);
   FAi_43 : FA_21 port map( A => A(43), B => B(43), Ci => tmp_43_port, S => 
                           S(43), Co => tmp_44_port);
   FAi_44 : FA_20 port map( A => A(44), B => B(44), Ci => tmp_44_port, S => 
                           S(44), Co => tmp_45_port);
   FAi_45 : FA_19 port map( A => A(45), B => B(45), Ci => tmp_45_port, S => 
                           S(45), Co => tmp_46_port);
   FAi_46 : FA_18 port map( A => A(46), B => B(46), Ci => tmp_46_port, S => 
                           S(46), Co => tmp_47_port);
   FAi_47 : FA_17 port map( A => A(47), B => B(47), Ci => tmp_47_port, S => 
                           S(47), Co => tmp_48_port);
   FAi_48 : FA_16 port map( A => A(48), B => B(48), Ci => tmp_48_port, S => 
                           S(48), Co => tmp_49_port);
   FAi_49 : FA_15 port map( A => A(49), B => B(49), Ci => tmp_49_port, S => 
                           S(49), Co => tmp_50_port);
   FAi_50 : FA_14 port map( A => A(50), B => B(50), Ci => tmp_50_port, S => 
                           S(50), Co => tmp_51_port);
   FAi_51 : FA_13 port map( A => A(51), B => B(51), Ci => tmp_51_port, S => 
                           S(51), Co => tmp_52_port);
   FAi_52 : FA_12 port map( A => A(52), B => B(52), Ci => tmp_52_port, S => 
                           S(52), Co => tmp_53_port);
   FAi_53 : FA_11 port map( A => A(53), B => B(53), Ci => tmp_53_port, S => 
                           S(53), Co => tmp_54_port);
   FAi_54 : FA_10 port map( A => A(54), B => B(54), Ci => tmp_54_port, S => 
                           S(54), Co => tmp_55_port);
   FAi_55 : FA_9 port map( A => A(55), B => B(55), Ci => tmp_55_port, S => 
                           S(55), Co => tmp_56_port);
   FAi_56 : FA_8 port map( A => A(56), B => B(56), Ci => tmp_56_port, S => 
                           S(56), Co => tmp_57_port);
   FAi_57 : FA_7 port map( A => A(57), B => B(57), Ci => tmp_57_port, S => 
                           S(57), Co => tmp_58_port);
   FAi_58 : FA_6 port map( A => A(58), B => B(58), Ci => tmp_58_port, S => 
                           S(58), Co => tmp_59_port);
   FAi_59 : FA_5 port map( A => A(59), B => B(59), Ci => tmp_59_port, S => 
                           S(59), Co => tmp_60_port);
   FAi_60 : FA_4 port map( A => A(60), B => B(60), Ci => tmp_60_port, S => 
                           S(60), Co => tmp_61_port);
   FAi_61 : FA_3 port map( A => A(61), B => B(61), Ci => tmp_61_port, S => 
                           S(61), Co => tmp_62_port);
   FAi_62 : FA_2 port map( A => A(62), B => B(62), Ci => tmp_62_port, S => 
                           S(62), Co => tmp_63_port);
   FAi_63 : FA_1 port map( A => A(63), B => B(63), Ci => tmp_63_port, S => 
                           S(63), Co => Co);

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity MUX21_GENERIC_N64 is

   port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y : 
         out std_logic_vector (63 downto 0));

end MUX21_GENERIC_N64;

architecture SYN_structural of MUX21_GENERIC_N64 is

   component NAND2_1
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_2
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_3
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_4
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_5
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_6
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_7
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_8
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_9
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_10
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_11
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_12
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_13
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_14
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_15
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_16
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_17
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_18
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_19
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_20
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_21
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_22
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_23
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_24
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_25
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_26
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_27
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_28
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_29
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_30
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_31
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_32
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_33
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_34
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_35
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_36
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_37
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_38
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_39
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_40
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_41
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_42
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_43
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_44
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_45
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_46
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_47
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_48
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_49
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_50
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_51
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_52
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_53
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_54
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_55
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_56
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_57
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_58
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_59
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_60
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_61
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_62
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_63
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_64
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_65
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_66
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_67
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_68
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_69
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_70
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_71
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_72
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_73
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_74
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_75
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_76
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_77
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_78
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_79
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_80
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_81
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_82
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_83
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_84
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_85
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_86
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_87
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_88
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_89
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_90
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_91
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_92
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_93
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_94
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_95
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_96
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_97
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_98
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_99
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_100
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_101
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_102
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_103
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_104
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_105
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_106
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_107
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_108
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_109
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_110
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_111
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_112
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_113
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_114
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_115
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_116
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_117
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_118
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_119
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_120
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_121
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_122
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_123
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_124
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_125
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_126
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_127
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_128
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_129
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_130
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_131
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_132
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_133
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_134
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_135
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_136
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_137
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_138
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_139
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_140
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_141
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_142
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_143
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_144
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_145
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_146
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_147
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_148
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_149
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_150
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_151
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_152
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_153
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_154
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_155
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_156
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_157
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_158
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_159
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_160
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_161
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_162
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_163
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_164
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_165
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_166
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_167
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_168
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_169
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_170
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_171
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_172
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_173
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_174
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_175
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_176
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_177
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_178
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_179
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_180
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_181
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_182
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_183
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_184
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_185
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_186
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_187
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_188
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_189
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_190
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_191
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component NAND2_0
      port( a, b : in std_logic;  f : out std_logic);
   end component;
   
   component INV
      port( a : in std_logic;  f : out std_logic);
   end component;
   
   signal sel_not, s1_63_port, s1_62_port, s1_61_port, s1_60_port, s1_59_port, 
      s1_58_port, s1_57_port, s1_56_port, s1_55_port, s1_54_port, s1_53_port, 
      s1_52_port, s1_51_port, s1_50_port, s1_49_port, s1_48_port, s1_47_port, 
      s1_46_port, s1_45_port, s1_44_port, s1_43_port, s1_42_port, s1_41_port, 
      s1_40_port, s1_39_port, s1_38_port, s1_37_port, s1_36_port, s1_35_port, 
      s1_34_port, s1_33_port, s1_32_port, s1_31_port, s1_30_port, s1_29_port, 
      s1_28_port, s1_27_port, s1_26_port, s1_25_port, s1_24_port, s1_23_port, 
      s1_22_port, s1_21_port, s1_20_port, s1_19_port, s1_18_port, s1_17_port, 
      s1_16_port, s1_15_port, s1_14_port, s1_13_port, s1_12_port, s1_11_port, 
      s1_10_port, s1_9_port, s1_8_port, s1_7_port, s1_6_port, s1_5_port, 
      s1_4_port, s1_3_port, s1_2_port, s1_1_port, s1_0_port, s2_63_port, 
      s2_62_port, s2_61_port, s2_60_port, s2_59_port, s2_58_port, s2_57_port, 
      s2_56_port, s2_55_port, s2_54_port, s2_53_port, s2_52_port, s2_51_port, 
      s2_50_port, s2_49_port, s2_48_port, s2_47_port, s2_46_port, s2_45_port, 
      s2_44_port, s2_43_port, s2_42_port, s2_41_port, s2_40_port, s2_39_port, 
      s2_38_port, s2_37_port, s2_36_port, s2_35_port, s2_34_port, s2_33_port, 
      s2_32_port, s2_31_port, s2_30_port, s2_29_port, s2_28_port, s2_27_port, 
      s2_26_port, s2_25_port, s2_24_port, s2_23_port, s2_22_port, s2_21_port, 
      s2_20_port, s2_19_port, s2_18_port, s2_17_port, s2_16_port, s2_15_port, 
      s2_14_port, s2_13_port, s2_12_port, s2_11_port, s2_10_port, s2_9_port, 
      s2_8_port, s2_7_port, s2_6_port, s2_5_port, s2_4_port, s2_3_port, 
      s2_2_port, s2_1_port, s2_0_port : std_logic;

begin
   
   inv_sel : INV port map( a => SEL, f => sel_not);
   s1_i_0 : NAND2_0 port map( a => A(0), b => sel_not, f => s1_0_port);
   s2_i_0 : NAND2_191 port map( a => B(0), b => SEL, f => s2_0_port);
   y_i_0 : NAND2_190 port map( a => s1_0_port, b => s2_0_port, f => Y(0));
   s1_i_1 : NAND2_189 port map( a => A(1), b => sel_not, f => s1_1_port);
   s2_i_1 : NAND2_188 port map( a => B(1), b => SEL, f => s2_1_port);
   y_i_1 : NAND2_187 port map( a => s1_1_port, b => s2_1_port, f => Y(1));
   s1_i_2 : NAND2_186 port map( a => A(2), b => sel_not, f => s1_2_port);
   s2_i_2 : NAND2_185 port map( a => B(2), b => SEL, f => s2_2_port);
   y_i_2 : NAND2_184 port map( a => s1_2_port, b => s2_2_port, f => Y(2));
   s1_i_3 : NAND2_183 port map( a => A(3), b => sel_not, f => s1_3_port);
   s2_i_3 : NAND2_182 port map( a => B(3), b => SEL, f => s2_3_port);
   y_i_3 : NAND2_181 port map( a => s1_3_port, b => s2_3_port, f => Y(3));
   s1_i_4 : NAND2_180 port map( a => A(4), b => sel_not, f => s1_4_port);
   s2_i_4 : NAND2_179 port map( a => B(4), b => SEL, f => s2_4_port);
   y_i_4 : NAND2_178 port map( a => s1_4_port, b => s2_4_port, f => Y(4));
   s1_i_5 : NAND2_177 port map( a => A(5), b => sel_not, f => s1_5_port);
   s2_i_5 : NAND2_176 port map( a => B(5), b => SEL, f => s2_5_port);
   y_i_5 : NAND2_175 port map( a => s1_5_port, b => s2_5_port, f => Y(5));
   s1_i_6 : NAND2_174 port map( a => A(6), b => sel_not, f => s1_6_port);
   s2_i_6 : NAND2_173 port map( a => B(6), b => SEL, f => s2_6_port);
   y_i_6 : NAND2_172 port map( a => s1_6_port, b => s2_6_port, f => Y(6));
   s1_i_7 : NAND2_171 port map( a => A(7), b => sel_not, f => s1_7_port);
   s2_i_7 : NAND2_170 port map( a => B(7), b => SEL, f => s2_7_port);
   y_i_7 : NAND2_169 port map( a => s1_7_port, b => s2_7_port, f => Y(7));
   s1_i_8 : NAND2_168 port map( a => A(8), b => sel_not, f => s1_8_port);
   s2_i_8 : NAND2_167 port map( a => B(8), b => SEL, f => s2_8_port);
   y_i_8 : NAND2_166 port map( a => s1_8_port, b => s2_8_port, f => Y(8));
   s1_i_9 : NAND2_165 port map( a => A(9), b => sel_not, f => s1_9_port);
   s2_i_9 : NAND2_164 port map( a => B(9), b => SEL, f => s2_9_port);
   y_i_9 : NAND2_163 port map( a => s1_9_port, b => s2_9_port, f => Y(9));
   s1_i_10 : NAND2_162 port map( a => A(10), b => sel_not, f => s1_10_port);
   s2_i_10 : NAND2_161 port map( a => B(10), b => SEL, f => s2_10_port);
   y_i_10 : NAND2_160 port map( a => s1_10_port, b => s2_10_port, f => Y(10));
   s1_i_11 : NAND2_159 port map( a => A(11), b => sel_not, f => s1_11_port);
   s2_i_11 : NAND2_158 port map( a => B(11), b => SEL, f => s2_11_port);
   y_i_11 : NAND2_157 port map( a => s1_11_port, b => s2_11_port, f => Y(11));
   s1_i_12 : NAND2_156 port map( a => A(12), b => sel_not, f => s1_12_port);
   s2_i_12 : NAND2_155 port map( a => B(12), b => SEL, f => s2_12_port);
   y_i_12 : NAND2_154 port map( a => s1_12_port, b => s2_12_port, f => Y(12));
   s1_i_13 : NAND2_153 port map( a => A(13), b => sel_not, f => s1_13_port);
   s2_i_13 : NAND2_152 port map( a => B(13), b => SEL, f => s2_13_port);
   y_i_13 : NAND2_151 port map( a => s1_13_port, b => s2_13_port, f => Y(13));
   s1_i_14 : NAND2_150 port map( a => A(14), b => sel_not, f => s1_14_port);
   s2_i_14 : NAND2_149 port map( a => B(14), b => SEL, f => s2_14_port);
   y_i_14 : NAND2_148 port map( a => s1_14_port, b => s2_14_port, f => Y(14));
   s1_i_15 : NAND2_147 port map( a => A(15), b => sel_not, f => s1_15_port);
   s2_i_15 : NAND2_146 port map( a => B(15), b => SEL, f => s2_15_port);
   y_i_15 : NAND2_145 port map( a => s1_15_port, b => s2_15_port, f => Y(15));
   s1_i_16 : NAND2_144 port map( a => A(16), b => sel_not, f => s1_16_port);
   s2_i_16 : NAND2_143 port map( a => B(16), b => SEL, f => s2_16_port);
   y_i_16 : NAND2_142 port map( a => s1_16_port, b => s2_16_port, f => Y(16));
   s1_i_17 : NAND2_141 port map( a => A(17), b => sel_not, f => s1_17_port);
   s2_i_17 : NAND2_140 port map( a => B(17), b => SEL, f => s2_17_port);
   y_i_17 : NAND2_139 port map( a => s1_17_port, b => s2_17_port, f => Y(17));
   s1_i_18 : NAND2_138 port map( a => A(18), b => sel_not, f => s1_18_port);
   s2_i_18 : NAND2_137 port map( a => B(18), b => SEL, f => s2_18_port);
   y_i_18 : NAND2_136 port map( a => s1_18_port, b => s2_18_port, f => Y(18));
   s1_i_19 : NAND2_135 port map( a => A(19), b => sel_not, f => s1_19_port);
   s2_i_19 : NAND2_134 port map( a => B(19), b => SEL, f => s2_19_port);
   y_i_19 : NAND2_133 port map( a => s1_19_port, b => s2_19_port, f => Y(19));
   s1_i_20 : NAND2_132 port map( a => A(20), b => sel_not, f => s1_20_port);
   s2_i_20 : NAND2_131 port map( a => B(20), b => SEL, f => s2_20_port);
   y_i_20 : NAND2_130 port map( a => s1_20_port, b => s2_20_port, f => Y(20));
   s1_i_21 : NAND2_129 port map( a => A(21), b => sel_not, f => s1_21_port);
   s2_i_21 : NAND2_128 port map( a => B(21), b => SEL, f => s2_21_port);
   y_i_21 : NAND2_127 port map( a => s1_21_port, b => s2_21_port, f => Y(21));
   s1_i_22 : NAND2_126 port map( a => A(22), b => sel_not, f => s1_22_port);
   s2_i_22 : NAND2_125 port map( a => B(22), b => SEL, f => s2_22_port);
   y_i_22 : NAND2_124 port map( a => s1_22_port, b => s2_22_port, f => Y(22));
   s1_i_23 : NAND2_123 port map( a => A(23), b => sel_not, f => s1_23_port);
   s2_i_23 : NAND2_122 port map( a => B(23), b => SEL, f => s2_23_port);
   y_i_23 : NAND2_121 port map( a => s1_23_port, b => s2_23_port, f => Y(23));
   s1_i_24 : NAND2_120 port map( a => A(24), b => sel_not, f => s1_24_port);
   s2_i_24 : NAND2_119 port map( a => B(24), b => SEL, f => s2_24_port);
   y_i_24 : NAND2_118 port map( a => s1_24_port, b => s2_24_port, f => Y(24));
   s1_i_25 : NAND2_117 port map( a => A(25), b => sel_not, f => s1_25_port);
   s2_i_25 : NAND2_116 port map( a => B(25), b => SEL, f => s2_25_port);
   y_i_25 : NAND2_115 port map( a => s1_25_port, b => s2_25_port, f => Y(25));
   s1_i_26 : NAND2_114 port map( a => A(26), b => sel_not, f => s1_26_port);
   s2_i_26 : NAND2_113 port map( a => B(26), b => SEL, f => s2_26_port);
   y_i_26 : NAND2_112 port map( a => s1_26_port, b => s2_26_port, f => Y(26));
   s1_i_27 : NAND2_111 port map( a => A(27), b => sel_not, f => s1_27_port);
   s2_i_27 : NAND2_110 port map( a => B(27), b => SEL, f => s2_27_port);
   y_i_27 : NAND2_109 port map( a => s1_27_port, b => s2_27_port, f => Y(27));
   s1_i_28 : NAND2_108 port map( a => A(28), b => sel_not, f => s1_28_port);
   s2_i_28 : NAND2_107 port map( a => B(28), b => SEL, f => s2_28_port);
   y_i_28 : NAND2_106 port map( a => s1_28_port, b => s2_28_port, f => Y(28));
   s1_i_29 : NAND2_105 port map( a => A(29), b => sel_not, f => s1_29_port);
   s2_i_29 : NAND2_104 port map( a => B(29), b => SEL, f => s2_29_port);
   y_i_29 : NAND2_103 port map( a => s1_29_port, b => s2_29_port, f => Y(29));
   s1_i_30 : NAND2_102 port map( a => A(30), b => sel_not, f => s1_30_port);
   s2_i_30 : NAND2_101 port map( a => B(30), b => SEL, f => s2_30_port);
   y_i_30 : NAND2_100 port map( a => s1_30_port, b => s2_30_port, f => Y(30));
   s1_i_31 : NAND2_99 port map( a => A(31), b => sel_not, f => s1_31_port);
   s2_i_31 : NAND2_98 port map( a => B(31), b => SEL, f => s2_31_port);
   y_i_31 : NAND2_97 port map( a => s1_31_port, b => s2_31_port, f => Y(31));
   s1_i_32 : NAND2_96 port map( a => A(32), b => sel_not, f => s1_32_port);
   s2_i_32 : NAND2_95 port map( a => B(32), b => SEL, f => s2_32_port);
   y_i_32 : NAND2_94 port map( a => s1_32_port, b => s2_32_port, f => Y(32));
   s1_i_33 : NAND2_93 port map( a => A(33), b => sel_not, f => s1_33_port);
   s2_i_33 : NAND2_92 port map( a => B(33), b => SEL, f => s2_33_port);
   y_i_33 : NAND2_91 port map( a => s1_33_port, b => s2_33_port, f => Y(33));
   s1_i_34 : NAND2_90 port map( a => A(34), b => sel_not, f => s1_34_port);
   s2_i_34 : NAND2_89 port map( a => B(34), b => SEL, f => s2_34_port);
   y_i_34 : NAND2_88 port map( a => s1_34_port, b => s2_34_port, f => Y(34));
   s1_i_35 : NAND2_87 port map( a => A(35), b => sel_not, f => s1_35_port);
   s2_i_35 : NAND2_86 port map( a => B(35), b => SEL, f => s2_35_port);
   y_i_35 : NAND2_85 port map( a => s1_35_port, b => s2_35_port, f => Y(35));
   s1_i_36 : NAND2_84 port map( a => A(36), b => sel_not, f => s1_36_port);
   s2_i_36 : NAND2_83 port map( a => B(36), b => SEL, f => s2_36_port);
   y_i_36 : NAND2_82 port map( a => s1_36_port, b => s2_36_port, f => Y(36));
   s1_i_37 : NAND2_81 port map( a => A(37), b => sel_not, f => s1_37_port);
   s2_i_37 : NAND2_80 port map( a => B(37), b => SEL, f => s2_37_port);
   y_i_37 : NAND2_79 port map( a => s1_37_port, b => s2_37_port, f => Y(37));
   s1_i_38 : NAND2_78 port map( a => A(38), b => sel_not, f => s1_38_port);
   s2_i_38 : NAND2_77 port map( a => B(38), b => SEL, f => s2_38_port);
   y_i_38 : NAND2_76 port map( a => s1_38_port, b => s2_38_port, f => Y(38));
   s1_i_39 : NAND2_75 port map( a => A(39), b => sel_not, f => s1_39_port);
   s2_i_39 : NAND2_74 port map( a => B(39), b => SEL, f => s2_39_port);
   y_i_39 : NAND2_73 port map( a => s1_39_port, b => s2_39_port, f => Y(39));
   s1_i_40 : NAND2_72 port map( a => A(40), b => sel_not, f => s1_40_port);
   s2_i_40 : NAND2_71 port map( a => B(40), b => SEL, f => s2_40_port);
   y_i_40 : NAND2_70 port map( a => s1_40_port, b => s2_40_port, f => Y(40));
   s1_i_41 : NAND2_69 port map( a => A(41), b => sel_not, f => s1_41_port);
   s2_i_41 : NAND2_68 port map( a => B(41), b => SEL, f => s2_41_port);
   y_i_41 : NAND2_67 port map( a => s1_41_port, b => s2_41_port, f => Y(41));
   s1_i_42 : NAND2_66 port map( a => A(42), b => sel_not, f => s1_42_port);
   s2_i_42 : NAND2_65 port map( a => B(42), b => SEL, f => s2_42_port);
   y_i_42 : NAND2_64 port map( a => s1_42_port, b => s2_42_port, f => Y(42));
   s1_i_43 : NAND2_63 port map( a => A(43), b => sel_not, f => s1_43_port);
   s2_i_43 : NAND2_62 port map( a => B(43), b => SEL, f => s2_43_port);
   y_i_43 : NAND2_61 port map( a => s1_43_port, b => s2_43_port, f => Y(43));
   s1_i_44 : NAND2_60 port map( a => A(44), b => sel_not, f => s1_44_port);
   s2_i_44 : NAND2_59 port map( a => B(44), b => SEL, f => s2_44_port);
   y_i_44 : NAND2_58 port map( a => s1_44_port, b => s2_44_port, f => Y(44));
   s1_i_45 : NAND2_57 port map( a => A(45), b => sel_not, f => s1_45_port);
   s2_i_45 : NAND2_56 port map( a => B(45), b => SEL, f => s2_45_port);
   y_i_45 : NAND2_55 port map( a => s1_45_port, b => s2_45_port, f => Y(45));
   s1_i_46 : NAND2_54 port map( a => A(46), b => sel_not, f => s1_46_port);
   s2_i_46 : NAND2_53 port map( a => B(46), b => SEL, f => s2_46_port);
   y_i_46 : NAND2_52 port map( a => s1_46_port, b => s2_46_port, f => Y(46));
   s1_i_47 : NAND2_51 port map( a => A(47), b => sel_not, f => s1_47_port);
   s2_i_47 : NAND2_50 port map( a => B(47), b => SEL, f => s2_47_port);
   y_i_47 : NAND2_49 port map( a => s1_47_port, b => s2_47_port, f => Y(47));
   s1_i_48 : NAND2_48 port map( a => A(48), b => sel_not, f => s1_48_port);
   s2_i_48 : NAND2_47 port map( a => B(48), b => SEL, f => s2_48_port);
   y_i_48 : NAND2_46 port map( a => s1_48_port, b => s2_48_port, f => Y(48));
   s1_i_49 : NAND2_45 port map( a => A(49), b => sel_not, f => s1_49_port);
   s2_i_49 : NAND2_44 port map( a => B(49), b => SEL, f => s2_49_port);
   y_i_49 : NAND2_43 port map( a => s1_49_port, b => s2_49_port, f => Y(49));
   s1_i_50 : NAND2_42 port map( a => A(50), b => sel_not, f => s1_50_port);
   s2_i_50 : NAND2_41 port map( a => B(50), b => SEL, f => s2_50_port);
   y_i_50 : NAND2_40 port map( a => s1_50_port, b => s2_50_port, f => Y(50));
   s1_i_51 : NAND2_39 port map( a => A(51), b => sel_not, f => s1_51_port);
   s2_i_51 : NAND2_38 port map( a => B(51), b => SEL, f => s2_51_port);
   y_i_51 : NAND2_37 port map( a => s1_51_port, b => s2_51_port, f => Y(51));
   s1_i_52 : NAND2_36 port map( a => A(52), b => sel_not, f => s1_52_port);
   s2_i_52 : NAND2_35 port map( a => B(52), b => SEL, f => s2_52_port);
   y_i_52 : NAND2_34 port map( a => s1_52_port, b => s2_52_port, f => Y(52));
   s1_i_53 : NAND2_33 port map( a => A(53), b => sel_not, f => s1_53_port);
   s2_i_53 : NAND2_32 port map( a => B(53), b => SEL, f => s2_53_port);
   y_i_53 : NAND2_31 port map( a => s1_53_port, b => s2_53_port, f => Y(53));
   s1_i_54 : NAND2_30 port map( a => A(54), b => sel_not, f => s1_54_port);
   s2_i_54 : NAND2_29 port map( a => B(54), b => SEL, f => s2_54_port);
   y_i_54 : NAND2_28 port map( a => s1_54_port, b => s2_54_port, f => Y(54));
   s1_i_55 : NAND2_27 port map( a => A(55), b => sel_not, f => s1_55_port);
   s2_i_55 : NAND2_26 port map( a => B(55), b => SEL, f => s2_55_port);
   y_i_55 : NAND2_25 port map( a => s1_55_port, b => s2_55_port, f => Y(55));
   s1_i_56 : NAND2_24 port map( a => A(56), b => sel_not, f => s1_56_port);
   s2_i_56 : NAND2_23 port map( a => B(56), b => SEL, f => s2_56_port);
   y_i_56 : NAND2_22 port map( a => s1_56_port, b => s2_56_port, f => Y(56));
   s1_i_57 : NAND2_21 port map( a => A(57), b => sel_not, f => s1_57_port);
   s2_i_57 : NAND2_20 port map( a => B(57), b => SEL, f => s2_57_port);
   y_i_57 : NAND2_19 port map( a => s1_57_port, b => s2_57_port, f => Y(57));
   s1_i_58 : NAND2_18 port map( a => A(58), b => sel_not, f => s1_58_port);
   s2_i_58 : NAND2_17 port map( a => B(58), b => SEL, f => s2_58_port);
   y_i_58 : NAND2_16 port map( a => s1_58_port, b => s2_58_port, f => Y(58));
   s1_i_59 : NAND2_15 port map( a => A(59), b => sel_not, f => s1_59_port);
   s2_i_59 : NAND2_14 port map( a => B(59), b => SEL, f => s2_59_port);
   y_i_59 : NAND2_13 port map( a => s1_59_port, b => s2_59_port, f => Y(59));
   s1_i_60 : NAND2_12 port map( a => A(60), b => sel_not, f => s1_60_port);
   s2_i_60 : NAND2_11 port map( a => B(60), b => SEL, f => s2_60_port);
   y_i_60 : NAND2_10 port map( a => s1_60_port, b => s2_60_port, f => Y(60));
   s1_i_61 : NAND2_9 port map( a => A(61), b => sel_not, f => s1_61_port);
   s2_i_61 : NAND2_8 port map( a => B(61), b => SEL, f => s2_61_port);
   y_i_61 : NAND2_7 port map( a => s1_61_port, b => s2_61_port, f => Y(61));
   s1_i_62 : NAND2_6 port map( a => A(62), b => sel_not, f => s1_62_port);
   s2_i_62 : NAND2_5 port map( a => B(62), b => SEL, f => s2_62_port);
   y_i_62 : NAND2_4 port map( a => s1_62_port, b => s2_62_port, f => Y(62));
   s1_i_63 : NAND2_3 port map( a => A(63), b => sel_not, f => s1_63_port);
   s2_i_63 : NAND2_2 port map( a => B(63), b => SEL, f => s2_63_port);
   y_i_63 : NAND2_1 port map( a => s1_63_port, b => s2_63_port, f => Y(63));

end SYN_structural;

library IEEE;

use IEEE.std_logic_1164.all;

use work.CONV_PACK_ACC_N64_1.all;

entity ACC_N64_1 is

   port( A, B : in std_logic_vector (63 downto 0);  CLK, RST_n, ACCUMULATE, 
         ACC_EN_n : in std_logic;  Y : out std_logic_vector (63 downto 0));

end ACC_N64_1;

architecture SYN_structural of ACC_N64_1 is

   component INV_X4
      port( A : in std_logic;  ZN : out std_logic);
   end component;
   
   component FD_GENERIC_N64
      port( D : in std_logic_vector (63 downto 0);  CK, RESET, ENABLE : in 
            std_logic;  Q : out std_logic_vector (63 downto 0));
   end component;
   
   component RCA_N64
      port( A, B : in std_logic_vector (63 downto 0);  Ci : in std_logic;  S : 
            out std_logic_vector (63 downto 0);  Co : out std_logic);
   end component;
   
   component MUX21_GENERIC_N64
      port( A, B : in std_logic_vector (63 downto 0);  SEL : in std_logic;  Y :
            out std_logic_vector (63 downto 0));
   end component;
   
   signal X_Logic0_port, Y_63_port, Y_62_port, Y_61_port, Y_60_port, Y_59_port,
      Y_58_port, Y_57_port, Y_56_port, Y_55_port, Y_54_port, Y_53_port, 
      Y_52_port, Y_51_port, Y_50_port, Y_49_port, Y_48_port, Y_47_port, 
      Y_46_port, Y_45_port, Y_44_port, Y_43_port, Y_42_port, Y_41_port, 
      Y_40_port, Y_39_port, Y_38_port, Y_37_port, Y_36_port, Y_35_port, 
      Y_34_port, Y_33_port, Y_32_port, Y_31_port, Y_30_port, Y_29_port, 
      Y_28_port, Y_27_port, Y_26_port, Y_25_port, Y_24_port, Y_23_port, 
      Y_22_port, Y_21_port, Y_20_port, Y_19_port, Y_18_port, Y_17_port, 
      Y_16_port, Y_15_port, Y_14_port, Y_13_port, Y_12_port, Y_11_port, 
      Y_10_port, Y_9_port, Y_8_port, Y_7_port, Y_6_port, Y_5_port, Y_4_port, 
      Y_3_port, Y_2_port, Y_1_port, Y_0_port, mux_out_63_port, mux_out_62_port,
      mux_out_61_port, mux_out_60_port, mux_out_59_port, mux_out_58_port, 
      mux_out_57_port, mux_out_56_port, mux_out_55_port, mux_out_54_port, 
      mux_out_53_port, mux_out_52_port, mux_out_51_port, mux_out_50_port, 
      mux_out_49_port, mux_out_48_port, mux_out_47_port, mux_out_46_port, 
      mux_out_45_port, mux_out_44_port, mux_out_43_port, mux_out_42_port, 
      mux_out_41_port, mux_out_40_port, mux_out_39_port, mux_out_38_port, 
      mux_out_37_port, mux_out_36_port, mux_out_35_port, mux_out_34_port, 
      mux_out_33_port, mux_out_32_port, mux_out_31_port, mux_out_30_port, 
      mux_out_29_port, mux_out_28_port, mux_out_27_port, mux_out_26_port, 
      mux_out_25_port, mux_out_24_port, mux_out_23_port, mux_out_22_port, 
      mux_out_21_port, mux_out_20_port, mux_out_19_port, mux_out_18_port, 
      mux_out_17_port, mux_out_16_port, mux_out_15_port, mux_out_14_port, 
      mux_out_13_port, mux_out_12_port, mux_out_11_port, mux_out_10_port, 
      mux_out_9_port, mux_out_8_port, mux_out_7_port, mux_out_6_port, 
      mux_out_5_port, mux_out_4_port, mux_out_3_port, mux_out_2_port, 
      mux_out_1_port, mux_out_0_port, out_add_63_port, out_add_62_port, 
      out_add_61_port, out_add_60_port, out_add_59_port, out_add_58_port, 
      out_add_57_port, out_add_56_port, out_add_55_port, out_add_54_port, 
      out_add_53_port, out_add_52_port, out_add_51_port, out_add_50_port, 
      out_add_49_port, out_add_48_port, out_add_47_port, out_add_46_port, 
      out_add_45_port, out_add_44_port, out_add_43_port, out_add_42_port, 
      out_add_41_port, out_add_40_port, out_add_39_port, out_add_38_port, 
      out_add_37_port, out_add_36_port, out_add_35_port, out_add_34_port, 
      out_add_33_port, out_add_32_port, out_add_31_port, out_add_30_port, 
      out_add_29_port, out_add_28_port, out_add_27_port, out_add_26_port, 
      out_add_25_port, out_add_24_port, out_add_23_port, out_add_22_port, 
      out_add_21_port, out_add_20_port, out_add_19_port, out_add_18_port, 
      out_add_17_port, out_add_16_port, out_add_15_port, out_add_14_port, 
      out_add_13_port, out_add_12_port, out_add_11_port, out_add_10_port, 
      out_add_9_port, out_add_8_port, out_add_7_port, out_add_6_port, 
      out_add_5_port, out_add_4_port, out_add_3_port, out_add_2_port, 
      out_add_1_port, out_add_0_port, n1, n2, n_1064 : std_logic;

begin
   Y <= ( Y_63_port, Y_62_port, Y_61_port, Y_60_port, Y_59_port, Y_58_port, 
      Y_57_port, Y_56_port, Y_55_port, Y_54_port, Y_53_port, Y_52_port, 
      Y_51_port, Y_50_port, Y_49_port, Y_48_port, Y_47_port, Y_46_port, 
      Y_45_port, Y_44_port, Y_43_port, Y_42_port, Y_41_port, Y_40_port, 
      Y_39_port, Y_38_port, Y_37_port, Y_36_port, Y_35_port, Y_34_port, 
      Y_33_port, Y_32_port, Y_31_port, Y_30_port, Y_29_port, Y_28_port, 
      Y_27_port, Y_26_port, Y_25_port, Y_24_port, Y_23_port, Y_22_port, 
      Y_21_port, Y_20_port, Y_19_port, Y_18_port, Y_17_port, Y_16_port, 
      Y_15_port, Y_14_port, Y_13_port, Y_12_port, Y_11_port, Y_10_port, 
      Y_9_port, Y_8_port, Y_7_port, Y_6_port, Y_5_port, Y_4_port, Y_3_port, 
      Y_2_port, Y_1_port, Y_0_port );
   
   mux : MUX21_GENERIC_N64 port map( A(63) => B(63), A(62) => B(62), A(61) => 
                           B(61), A(60) => B(60), A(59) => B(59), A(58) => 
                           B(58), A(57) => B(57), A(56) => B(56), A(55) => 
                           B(55), A(54) => B(54), A(53) => B(53), A(52) => 
                           B(52), A(51) => B(51), A(50) => B(50), A(49) => 
                           B(49), A(48) => B(48), A(47) => B(47), A(46) => 
                           B(46), A(45) => B(45), A(44) => B(44), A(43) => 
                           B(43), A(42) => B(42), A(41) => B(41), A(40) => 
                           B(40), A(39) => B(39), A(38) => B(38), A(37) => 
                           B(37), A(36) => B(36), A(35) => B(35), A(34) => 
                           B(34), A(33) => B(33), A(32) => B(32), A(31) => 
                           B(31), A(30) => B(30), A(29) => B(29), A(28) => 
                           B(28), A(27) => B(27), A(26) => B(26), A(25) => 
                           B(25), A(24) => B(24), A(23) => B(23), A(22) => 
                           B(22), A(21) => B(21), A(20) => B(20), A(19) => 
                           B(19), A(18) => B(18), A(17) => B(17), A(16) => 
                           B(16), A(15) => B(15), A(14) => B(14), A(13) => 
                           B(13), A(12) => B(12), A(11) => B(11), A(10) => 
                           B(10), A(9) => B(9), A(8) => B(8), A(7) => B(7), 
                           A(6) => B(6), A(5) => B(5), A(4) => B(4), A(3) => 
                           B(3), A(2) => B(2), A(1) => B(1), A(0) => B(0), 
                           B(63) => Y_63_port, B(62) => Y_62_port, B(61) => 
                           Y_61_port, B(60) => Y_60_port, B(59) => Y_59_port, 
                           B(58) => Y_58_port, B(57) => Y_57_port, B(56) => 
                           Y_56_port, B(55) => Y_55_port, B(54) => Y_54_port, 
                           B(53) => Y_53_port, B(52) => Y_52_port, B(51) => 
                           Y_51_port, B(50) => Y_50_port, B(49) => Y_49_port, 
                           B(48) => Y_48_port, B(47) => Y_47_port, B(46) => 
                           Y_46_port, B(45) => Y_45_port, B(44) => Y_44_port, 
                           B(43) => Y_43_port, B(42) => Y_42_port, B(41) => 
                           Y_41_port, B(40) => Y_40_port, B(39) => Y_39_port, 
                           B(38) => Y_38_port, B(37) => Y_37_port, B(36) => 
                           Y_36_port, B(35) => Y_35_port, B(34) => Y_34_port, 
                           B(33) => Y_33_port, B(32) => Y_32_port, B(31) => 
                           Y_31_port, B(30) => Y_30_port, B(29) => Y_29_port, 
                           B(28) => Y_28_port, B(27) => Y_27_port, B(26) => 
                           Y_26_port, B(25) => Y_25_port, B(24) => Y_24_port, 
                           B(23) => Y_23_port, B(22) => Y_22_port, B(21) => 
                           Y_21_port, B(20) => Y_20_port, B(19) => Y_19_port, 
                           B(18) => Y_18_port, B(17) => Y_17_port, B(16) => 
                           Y_16_port, B(15) => Y_15_port, B(14) => Y_14_port, 
                           B(13) => Y_13_port, B(12) => Y_12_port, B(11) => 
                           Y_11_port, B(10) => Y_10_port, B(9) => Y_9_port, 
                           B(8) => Y_8_port, B(7) => Y_7_port, B(6) => Y_6_port
                           , B(5) => Y_5_port, B(4) => Y_4_port, B(3) => 
                           Y_3_port, B(2) => Y_2_port, B(1) => Y_1_port, B(0) 
                           => Y_0_port, SEL => ACCUMULATE, Y(63) => 
                           mux_out_63_port, Y(62) => mux_out_62_port, Y(61) => 
                           mux_out_61_port, Y(60) => mux_out_60_port, Y(59) => 
                           mux_out_59_port, Y(58) => mux_out_58_port, Y(57) => 
                           mux_out_57_port, Y(56) => mux_out_56_port, Y(55) => 
                           mux_out_55_port, Y(54) => mux_out_54_port, Y(53) => 
                           mux_out_53_port, Y(52) => mux_out_52_port, Y(51) => 
                           mux_out_51_port, Y(50) => mux_out_50_port, Y(49) => 
                           mux_out_49_port, Y(48) => mux_out_48_port, Y(47) => 
                           mux_out_47_port, Y(46) => mux_out_46_port, Y(45) => 
                           mux_out_45_port, Y(44) => mux_out_44_port, Y(43) => 
                           mux_out_43_port, Y(42) => mux_out_42_port, Y(41) => 
                           mux_out_41_port, Y(40) => mux_out_40_port, Y(39) => 
                           mux_out_39_port, Y(38) => mux_out_38_port, Y(37) => 
                           mux_out_37_port, Y(36) => mux_out_36_port, Y(35) => 
                           mux_out_35_port, Y(34) => mux_out_34_port, Y(33) => 
                           mux_out_33_port, Y(32) => mux_out_32_port, Y(31) => 
                           mux_out_31_port, Y(30) => mux_out_30_port, Y(29) => 
                           mux_out_29_port, Y(28) => mux_out_28_port, Y(27) => 
                           mux_out_27_port, Y(26) => mux_out_26_port, Y(25) => 
                           mux_out_25_port, Y(24) => mux_out_24_port, Y(23) => 
                           mux_out_23_port, Y(22) => mux_out_22_port, Y(21) => 
                           mux_out_21_port, Y(20) => mux_out_20_port, Y(19) => 
                           mux_out_19_port, Y(18) => mux_out_18_port, Y(17) => 
                           mux_out_17_port, Y(16) => mux_out_16_port, Y(15) => 
                           mux_out_15_port, Y(14) => mux_out_14_port, Y(13) => 
                           mux_out_13_port, Y(12) => mux_out_12_port, Y(11) => 
                           mux_out_11_port, Y(10) => mux_out_10_port, Y(9) => 
                           mux_out_9_port, Y(8) => mux_out_8_port, Y(7) => 
                           mux_out_7_port, Y(6) => mux_out_6_port, Y(5) => 
                           mux_out_5_port, Y(4) => mux_out_4_port, Y(3) => 
                           mux_out_3_port, Y(2) => mux_out_2_port, Y(1) => 
                           mux_out_1_port, Y(0) => mux_out_0_port);
   add : RCA_N64 port map( A(63) => A(63), A(62) => A(62), A(61) => A(61), 
                           A(60) => A(60), A(59) => A(59), A(58) => A(58), 
                           A(57) => A(57), A(56) => A(56), A(55) => A(55), 
                           A(54) => A(54), A(53) => A(53), A(52) => A(52), 
                           A(51) => A(51), A(50) => A(50), A(49) => A(49), 
                           A(48) => A(48), A(47) => A(47), A(46) => A(46), 
                           A(45) => A(45), A(44) => A(44), A(43) => A(43), 
                           A(42) => A(42), A(41) => A(41), A(40) => A(40), 
                           A(39) => A(39), A(38) => A(38), A(37) => A(37), 
                           A(36) => A(36), A(35) => A(35), A(34) => A(34), 
                           A(33) => A(33), A(32) => A(32), A(31) => A(31), 
                           A(30) => A(30), A(29) => A(29), A(28) => A(28), 
                           A(27) => A(27), A(26) => A(26), A(25) => A(25), 
                           A(24) => A(24), A(23) => A(23), A(22) => A(22), 
                           A(21) => A(21), A(20) => A(20), A(19) => A(19), 
                           A(18) => A(18), A(17) => A(17), A(16) => A(16), 
                           A(15) => A(15), A(14) => A(14), A(13) => A(13), 
                           A(12) => A(12), A(11) => A(11), A(10) => A(10), A(9)
                           => A(9), A(8) => A(8), A(7) => A(7), A(6) => A(6), 
                           A(5) => A(5), A(4) => A(4), A(3) => A(3), A(2) => 
                           A(2), A(1) => A(1), A(0) => A(0), B(63) => 
                           mux_out_63_port, B(62) => mux_out_62_port, B(61) => 
                           mux_out_61_port, B(60) => mux_out_60_port, B(59) => 
                           mux_out_59_port, B(58) => mux_out_58_port, B(57) => 
                           mux_out_57_port, B(56) => mux_out_56_port, B(55) => 
                           mux_out_55_port, B(54) => mux_out_54_port, B(53) => 
                           mux_out_53_port, B(52) => mux_out_52_port, B(51) => 
                           mux_out_51_port, B(50) => mux_out_50_port, B(49) => 
                           mux_out_49_port, B(48) => mux_out_48_port, B(47) => 
                           mux_out_47_port, B(46) => mux_out_46_port, B(45) => 
                           mux_out_45_port, B(44) => mux_out_44_port, B(43) => 
                           mux_out_43_port, B(42) => mux_out_42_port, B(41) => 
                           mux_out_41_port, B(40) => mux_out_40_port, B(39) => 
                           mux_out_39_port, B(38) => mux_out_38_port, B(37) => 
                           mux_out_37_port, B(36) => mux_out_36_port, B(35) => 
                           mux_out_35_port, B(34) => mux_out_34_port, B(33) => 
                           mux_out_33_port, B(32) => mux_out_32_port, B(31) => 
                           mux_out_31_port, B(30) => mux_out_30_port, B(29) => 
                           mux_out_29_port, B(28) => mux_out_28_port, B(27) => 
                           mux_out_27_port, B(26) => mux_out_26_port, B(25) => 
                           mux_out_25_port, B(24) => mux_out_24_port, B(23) => 
                           mux_out_23_port, B(22) => mux_out_22_port, B(21) => 
                           mux_out_21_port, B(20) => mux_out_20_port, B(19) => 
                           mux_out_19_port, B(18) => mux_out_18_port, B(17) => 
                           mux_out_17_port, B(16) => mux_out_16_port, B(15) => 
                           mux_out_15_port, B(14) => mux_out_14_port, B(13) => 
                           mux_out_13_port, B(12) => mux_out_12_port, B(11) => 
                           mux_out_11_port, B(10) => mux_out_10_port, B(9) => 
                           mux_out_9_port, B(8) => mux_out_8_port, B(7) => 
                           mux_out_7_port, B(6) => mux_out_6_port, B(5) => 
                           mux_out_5_port, B(4) => mux_out_4_port, B(3) => 
                           mux_out_3_port, B(2) => mux_out_2_port, B(1) => 
                           mux_out_1_port, B(0) => mux_out_0_port, Ci => 
                           X_Logic0_port, S(63) => out_add_63_port, S(62) => 
                           out_add_62_port, S(61) => out_add_61_port, S(60) => 
                           out_add_60_port, S(59) => out_add_59_port, S(58) => 
                           out_add_58_port, S(57) => out_add_57_port, S(56) => 
                           out_add_56_port, S(55) => out_add_55_port, S(54) => 
                           out_add_54_port, S(53) => out_add_53_port, S(52) => 
                           out_add_52_port, S(51) => out_add_51_port, S(50) => 
                           out_add_50_port, S(49) => out_add_49_port, S(48) => 
                           out_add_48_port, S(47) => out_add_47_port, S(46) => 
                           out_add_46_port, S(45) => out_add_45_port, S(44) => 
                           out_add_44_port, S(43) => out_add_43_port, S(42) => 
                           out_add_42_port, S(41) => out_add_41_port, S(40) => 
                           out_add_40_port, S(39) => out_add_39_port, S(38) => 
                           out_add_38_port, S(37) => out_add_37_port, S(36) => 
                           out_add_36_port, S(35) => out_add_35_port, S(34) => 
                           out_add_34_port, S(33) => out_add_33_port, S(32) => 
                           out_add_32_port, S(31) => out_add_31_port, S(30) => 
                           out_add_30_port, S(29) => out_add_29_port, S(28) => 
                           out_add_28_port, S(27) => out_add_27_port, S(26) => 
                           out_add_26_port, S(25) => out_add_25_port, S(24) => 
                           out_add_24_port, S(23) => out_add_23_port, S(22) => 
                           out_add_22_port, S(21) => out_add_21_port, S(20) => 
                           out_add_20_port, S(19) => out_add_19_port, S(18) => 
                           out_add_18_port, S(17) => out_add_17_port, S(16) => 
                           out_add_16_port, S(15) => out_add_15_port, S(14) => 
                           out_add_14_port, S(13) => out_add_13_port, S(12) => 
                           out_add_12_port, S(11) => out_add_11_port, S(10) => 
                           out_add_10_port, S(9) => out_add_9_port, S(8) => 
                           out_add_8_port, S(7) => out_add_7_port, S(6) => 
                           out_add_6_port, S(5) => out_add_5_port, S(4) => 
                           out_add_4_port, S(3) => out_add_3_port, S(2) => 
                           out_add_2_port, S(1) => out_add_1_port, S(0) => 
                           out_add_0_port, Co => n_1064);
   reg : FD_GENERIC_N64 port map( D(63) => out_add_63_port, D(62) => 
                           out_add_62_port, D(61) => out_add_61_port, D(60) => 
                           out_add_60_port, D(59) => out_add_59_port, D(58) => 
                           out_add_58_port, D(57) => out_add_57_port, D(56) => 
                           out_add_56_port, D(55) => out_add_55_port, D(54) => 
                           out_add_54_port, D(53) => out_add_53_port, D(52) => 
                           out_add_52_port, D(51) => out_add_51_port, D(50) => 
                           out_add_50_port, D(49) => out_add_49_port, D(48) => 
                           out_add_48_port, D(47) => out_add_47_port, D(46) => 
                           out_add_46_port, D(45) => out_add_45_port, D(44) => 
                           out_add_44_port, D(43) => out_add_43_port, D(42) => 
                           out_add_42_port, D(41) => out_add_41_port, D(40) => 
                           out_add_40_port, D(39) => out_add_39_port, D(38) => 
                           out_add_38_port, D(37) => out_add_37_port, D(36) => 
                           out_add_36_port, D(35) => out_add_35_port, D(34) => 
                           out_add_34_port, D(33) => out_add_33_port, D(32) => 
                           out_add_32_port, D(31) => out_add_31_port, D(30) => 
                           out_add_30_port, D(29) => out_add_29_port, D(28) => 
                           out_add_28_port, D(27) => out_add_27_port, D(26) => 
                           out_add_26_port, D(25) => out_add_25_port, D(24) => 
                           out_add_24_port, D(23) => out_add_23_port, D(22) => 
                           out_add_22_port, D(21) => out_add_21_port, D(20) => 
                           out_add_20_port, D(19) => out_add_19_port, D(18) => 
                           out_add_18_port, D(17) => out_add_17_port, D(16) => 
                           out_add_16_port, D(15) => out_add_15_port, D(14) => 
                           out_add_14_port, D(13) => out_add_13_port, D(12) => 
                           out_add_12_port, D(11) => out_add_11_port, D(10) => 
                           out_add_10_port, D(9) => out_add_9_port, D(8) => 
                           out_add_8_port, D(7) => out_add_7_port, D(6) => 
                           out_add_6_port, D(5) => out_add_5_port, D(4) => 
                           out_add_4_port, D(3) => out_add_3_port, D(2) => 
                           out_add_2_port, D(1) => out_add_1_port, D(0) => 
                           out_add_0_port, CK => CLK, RESET => n1, ENABLE => n2
                           , Q(63) => Y_63_port, Q(62) => Y_62_port, Q(61) => 
                           Y_61_port, Q(60) => Y_60_port, Q(59) => Y_59_port, 
                           Q(58) => Y_58_port, Q(57) => Y_57_port, Q(56) => 
                           Y_56_port, Q(55) => Y_55_port, Q(54) => Y_54_port, 
                           Q(53) => Y_53_port, Q(52) => Y_52_port, Q(51) => 
                           Y_51_port, Q(50) => Y_50_port, Q(49) => Y_49_port, 
                           Q(48) => Y_48_port, Q(47) => Y_47_port, Q(46) => 
                           Y_46_port, Q(45) => Y_45_port, Q(44) => Y_44_port, 
                           Q(43) => Y_43_port, Q(42) => Y_42_port, Q(41) => 
                           Y_41_port, Q(40) => Y_40_port, Q(39) => Y_39_port, 
                           Q(38) => Y_38_port, Q(37) => Y_37_port, Q(36) => 
                           Y_36_port, Q(35) => Y_35_port, Q(34) => Y_34_port, 
                           Q(33) => Y_33_port, Q(32) => Y_32_port, Q(31) => 
                           Y_31_port, Q(30) => Y_30_port, Q(29) => Y_29_port, 
                           Q(28) => Y_28_port, Q(27) => Y_27_port, Q(26) => 
                           Y_26_port, Q(25) => Y_25_port, Q(24) => Y_24_port, 
                           Q(23) => Y_23_port, Q(22) => Y_22_port, Q(21) => 
                           Y_21_port, Q(20) => Y_20_port, Q(19) => Y_19_port, 
                           Q(18) => Y_18_port, Q(17) => Y_17_port, Q(16) => 
                           Y_16_port, Q(15) => Y_15_port, Q(14) => Y_14_port, 
                           Q(13) => Y_13_port, Q(12) => Y_12_port, Q(11) => 
                           Y_11_port, Q(10) => Y_10_port, Q(9) => Y_9_port, 
                           Q(8) => Y_8_port, Q(7) => Y_7_port, Q(6) => Y_6_port
                           , Q(5) => Y_5_port, Q(4) => Y_4_port, Q(3) => 
                           Y_3_port, Q(2) => Y_2_port, Q(1) => Y_1_port, Q(0) 
                           => Y_0_port);
   X_Logic0_port <= '0';
   U4 : INV_X4 port map( A => RST_n, ZN => n1);
   U5 : INV_X4 port map( A => ACC_EN_n, ZN => n2);

end SYN_structural;
