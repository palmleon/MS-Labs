package CONSTANTS is
   -- kept  only used constants
   constant NumBit : integer := 4;	
   constant RAD : integer := 3;	
end CONSTANTS;
