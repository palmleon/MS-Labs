library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;
use IEEE.math_real.all;
use WORK.constants.all;

entity ThermometricDecoder32 is
    port 
    (
        IN1 : in std_logic_vector(4 downto 0);
        OUT1 : out std_logic_vector(31 downto 0)
    );
end entity;

architecture behavioral of ThermometricDecoder32 is
    begin
        process (IN1) 
        begin
            case IN1 is
                when "00000" => OUT1 <= "00000000000000000000000000000000";
                when "00001" => OUT1 <= "00000000000000000000000000000001";
                when "00010" => OUT1 <= "00000000000000000000000000000011";
                when "00011" => OUT1 <= "00000000000000000000000000000111";
                when "00100" => OUT1 <= "00000000000000000000000000001111";
                when "00101" => OUT1 <= "00000000000000000000000000011111";
                when "00110" => OUT1 <= "00000000000000000000000000111111";
                when "00111" => OUT1 <= "00000000000000000000000001111111";
                when "01000" => OUT1 <= "00000000000000000000000011111111";
                when "01001" => OUT1 <= "00000000000000000000000111111111";
                when "01010" => OUT1 <= "00000000000000000000001111111111";
                when "01011" => OUT1 <= "00000000000000000000011111111111";
                when "01100" => OUT1 <= "00000000000000000000111111111111";
                when "01101" => OUT1 <= "00000000000000000001111111111111";
                when "01110" => OUT1 <= "00000000000000000011111111111111";
                when "01111" => OUT1 <= "00000000000000000111111111111111";
                when "10000" => OUT1 <= "00000000000000001111111111111111";
                when "10001" => OUT1 <= "00000000000000011111111111111111";
                when "10010" => OUT1 <= "00000000000000111111111111111111";
                when "10011" => OUT1 <= "00000000000001111111111111111111";
                when "10100" => OUT1 <= "00000000000011111111111111111111";
                when "10101" => OUT1 <= "00000000000111111111111111111111";
                when "10110" => OUT1 <= "00000000001111111111111111111111";
                when "10111" => OUT1 <= "00000000011111111111111111111111";
                when "11000" => OUT1 <= "00000000111111111111111111111111";
                when "11001" => OUT1 <= "00000001111111111111111111111111";
                when "11010" => OUT1 <= "00000011111111111111111111111111";
                when "11011" => OUT1 <= "00000111111111111111111111111111";
                when "11100" => OUT1 <= "00001111111111111111111111111111";
                when "11101" => OUT1 <= "00011111111111111111111111111111";
                when "11110" => OUT1 <= "00111111111111111111111111111111";
                when "11111" => OUT1 <= "01111111111111111111111111111111";
                when others => OUT1 <= (others => '0');
            end case;
        end process;

end architecture;